magic
tech scmos
timestamp 1523021392
<< pwell >>
rect 495 230 543 256
rect 722 232 826 258
rect 855 232 903 258
rect 356 194 474 230
rect 36 89 179 114
rect 18 78 179 89
rect 486 194 629 230
rect 716 196 834 232
rect 846 196 989 232
rect 191 78 309 114
rect 392 104 526 106
rect 542 104 665 106
rect 392 82 665 104
rect 18 53 170 78
rect 392 70 535 82
rect 547 70 665 82
rect 752 106 886 108
rect 902 106 1025 108
rect 752 84 1025 106
rect 752 72 895 84
rect 907 72 1025 84
rect 122 52 170 53
rect 478 44 526 70
rect 838 46 886 72
<< nwell >>
rect 495 276 543 299
rect 495 263 547 276
rect 495 256 543 263
rect 722 258 826 302
rect 855 278 903 301
rect 855 265 907 278
rect 855 258 903 265
rect 36 114 179 158
rect 191 114 309 158
rect 356 154 474 194
rect 486 157 629 194
rect 486 154 664 157
rect 356 150 664 154
rect 716 156 834 196
rect 846 159 989 196
rect 846 156 1024 159
rect 716 152 1024 156
rect 358 145 665 150
rect 718 147 1025 152
rect 392 106 665 145
rect 526 104 542 106
rect 752 108 1025 147
rect 886 106 902 108
rect 18 52 122 53
rect 18 9 170 52
rect 478 37 526 44
rect 838 39 886 46
rect 474 24 526 37
rect 834 26 886 39
rect 122 8 170 9
rect 478 0 526 24
rect 838 2 886 26
<< polysilicon >>
rect 521 290 523 294
rect 528 290 530 294
rect 735 292 737 296
rect 508 281 510 285
rect 508 260 510 269
rect 521 267 523 272
rect 518 266 524 267
rect 518 262 519 266
rect 523 262 524 266
rect 518 261 524 262
rect 508 259 514 260
rect 508 255 509 259
rect 513 255 514 259
rect 518 258 520 261
rect 528 259 530 272
rect 758 289 760 309
rect 765 289 767 294
rect 783 292 785 296
rect 793 292 795 296
rect 803 292 805 296
rect 748 280 750 285
rect 528 258 534 259
rect 508 254 514 255
rect 528 254 529 258
rect 533 254 534 258
rect 508 245 510 254
rect 518 245 520 254
rect 528 253 534 254
rect 735 254 737 267
rect 748 264 750 267
rect 881 292 883 296
rect 888 292 890 296
rect 868 283 870 287
rect 741 263 750 264
rect 741 259 742 263
rect 746 262 750 263
rect 746 259 747 262
rect 758 261 760 264
rect 741 258 747 259
rect 735 253 741 254
rect 528 245 530 253
rect 735 249 736 253
rect 740 249 741 253
rect 735 248 741 249
rect 735 245 737 248
rect 745 245 747 258
rect 755 260 760 261
rect 755 256 756 260
rect 755 255 760 256
rect 765 261 767 264
rect 783 261 785 264
rect 793 261 795 264
rect 803 261 805 264
rect 868 262 870 271
rect 881 269 883 274
rect 878 268 884 269
rect 878 264 879 268
rect 883 264 884 268
rect 878 263 884 264
rect 868 261 874 262
rect 765 260 787 261
rect 765 256 775 260
rect 779 256 782 260
rect 786 256 787 260
rect 765 255 787 256
rect 791 260 797 261
rect 791 256 792 260
rect 796 256 797 260
rect 791 255 797 256
rect 801 260 807 261
rect 801 256 802 260
rect 806 256 807 260
rect 801 255 807 256
rect 868 257 869 261
rect 873 257 874 261
rect 878 260 880 263
rect 888 261 890 274
rect 888 260 894 261
rect 868 256 874 257
rect 888 256 889 260
rect 893 256 894 260
rect 755 252 757 255
rect 765 252 767 255
rect 785 252 787 255
rect 792 252 794 255
rect 508 235 510 239
rect 518 235 520 239
rect 528 235 530 239
rect 735 228 737 232
rect 745 230 747 235
rect 755 233 757 238
rect 765 233 767 238
rect 803 246 805 255
rect 868 247 870 256
rect 878 247 880 256
rect 888 255 894 256
rect 888 247 890 255
rect 868 237 870 241
rect 878 237 880 241
rect 888 237 890 241
rect 785 228 787 232
rect 792 228 794 232
rect 803 228 805 232
rect 370 217 372 222
rect 377 217 379 222
rect 433 222 458 224
rect 416 217 418 222
rect 423 217 425 222
rect 389 211 391 215
rect 370 205 372 208
rect 366 204 372 205
rect 366 200 367 204
rect 371 200 372 204
rect 366 199 372 200
rect 369 188 371 199
rect 377 194 379 208
rect 433 214 435 222
rect 443 214 445 218
rect 456 214 458 222
rect 517 222 542 224
rect 500 217 502 222
rect 507 217 509 222
rect 456 212 461 214
rect 459 209 461 212
rect 389 197 391 205
rect 385 196 391 197
rect 416 196 418 205
rect 423 202 425 205
rect 423 200 427 202
rect 433 200 435 205
rect 443 202 445 205
rect 443 201 452 202
rect 425 196 427 200
rect 443 197 447 201
rect 451 197 452 201
rect 517 214 519 222
rect 527 214 529 218
rect 540 214 542 222
rect 602 217 604 222
rect 609 217 611 222
rect 730 219 732 224
rect 737 219 739 224
rect 793 224 818 226
rect 776 219 778 224
rect 783 219 785 224
rect 540 212 545 214
rect 543 209 545 212
rect 443 196 452 197
rect 377 191 381 194
rect 385 192 386 196
rect 390 192 391 196
rect 385 191 391 192
rect 379 188 381 191
rect 389 188 391 191
rect 415 195 421 196
rect 415 191 416 195
rect 420 191 421 195
rect 415 190 421 191
rect 425 195 431 196
rect 425 191 426 195
rect 430 191 431 195
rect 443 192 445 196
rect 459 192 461 200
rect 500 196 502 205
rect 507 202 509 205
rect 507 200 511 202
rect 517 200 519 205
rect 527 202 529 205
rect 527 201 536 202
rect 509 196 511 200
rect 527 197 531 201
rect 535 197 536 201
rect 621 211 623 215
rect 602 205 604 208
rect 598 204 604 205
rect 598 200 599 204
rect 603 200 604 204
rect 527 196 536 197
rect 499 195 505 196
rect 425 190 431 191
rect 435 190 445 192
rect 451 190 464 192
rect 369 173 371 178
rect 379 173 381 178
rect 415 187 417 190
rect 425 187 427 190
rect 435 187 437 190
rect 451 187 453 190
rect 375 172 381 173
rect 375 168 376 172
rect 380 168 381 172
rect 389 171 391 176
rect 375 167 381 168
rect 425 165 427 169
rect 435 165 437 169
rect 415 156 417 160
rect 462 181 464 190
rect 499 191 500 195
rect 504 191 505 195
rect 499 190 505 191
rect 509 195 515 196
rect 509 191 510 195
rect 514 191 515 195
rect 527 192 529 196
rect 543 192 545 200
rect 598 199 604 200
rect 509 190 515 191
rect 519 190 529 192
rect 535 190 548 192
rect 499 187 501 190
rect 509 187 511 190
rect 519 187 521 190
rect 535 187 537 190
rect 462 180 468 181
rect 462 176 463 180
rect 467 176 468 180
rect 462 175 468 176
rect 509 165 511 169
rect 519 165 521 169
rect 451 156 453 160
rect 499 156 501 160
rect 546 181 548 190
rect 601 188 603 199
rect 609 194 611 208
rect 749 213 751 217
rect 730 207 732 210
rect 726 206 732 207
rect 621 197 623 205
rect 726 202 727 206
rect 731 202 732 206
rect 726 201 732 202
rect 617 196 623 197
rect 609 191 613 194
rect 617 192 618 196
rect 622 192 623 196
rect 617 191 623 192
rect 611 188 613 191
rect 621 188 623 191
rect 729 190 731 201
rect 737 196 739 210
rect 793 216 795 224
rect 803 216 805 220
rect 816 216 818 224
rect 877 224 902 226
rect 860 219 862 224
rect 867 219 869 224
rect 816 214 821 216
rect 819 211 821 214
rect 749 199 751 207
rect 745 198 751 199
rect 776 198 778 207
rect 783 204 785 207
rect 783 202 787 204
rect 793 202 795 207
rect 803 204 805 207
rect 803 203 812 204
rect 785 198 787 202
rect 803 199 807 203
rect 811 199 812 203
rect 877 216 879 224
rect 887 216 889 220
rect 900 216 902 224
rect 962 219 964 224
rect 969 219 971 224
rect 900 214 905 216
rect 903 211 905 214
rect 803 198 812 199
rect 737 193 741 196
rect 745 194 746 198
rect 750 194 751 198
rect 745 193 751 194
rect 739 190 741 193
rect 749 190 751 193
rect 775 197 781 198
rect 775 193 776 197
rect 780 193 781 197
rect 775 192 781 193
rect 785 197 791 198
rect 785 193 786 197
rect 790 193 791 197
rect 803 194 805 198
rect 819 194 821 202
rect 860 198 862 207
rect 867 204 869 207
rect 867 202 871 204
rect 877 202 879 207
rect 887 204 889 207
rect 887 203 896 204
rect 869 198 871 202
rect 887 199 891 203
rect 895 199 896 203
rect 981 213 983 217
rect 962 207 964 210
rect 958 206 964 207
rect 958 202 959 206
rect 963 202 964 206
rect 887 198 896 199
rect 859 197 865 198
rect 785 192 791 193
rect 795 192 805 194
rect 811 192 824 194
rect 546 180 552 181
rect 546 176 547 180
rect 551 176 552 180
rect 546 175 552 176
rect 601 173 603 178
rect 611 173 613 178
rect 607 172 613 173
rect 607 168 608 172
rect 612 168 613 172
rect 621 171 623 176
rect 729 175 731 180
rect 739 175 741 180
rect 775 189 777 192
rect 785 189 787 192
rect 795 189 797 192
rect 811 189 813 192
rect 735 174 741 175
rect 735 170 736 174
rect 740 170 741 174
rect 749 173 751 178
rect 735 169 741 170
rect 607 167 613 168
rect 535 156 537 160
rect 785 167 787 171
rect 795 167 797 171
rect 775 158 777 162
rect 822 183 824 192
rect 859 193 860 197
rect 864 193 865 197
rect 859 192 865 193
rect 869 197 875 198
rect 869 193 870 197
rect 874 193 875 197
rect 887 194 889 198
rect 903 194 905 202
rect 958 201 964 202
rect 869 192 875 193
rect 879 192 889 194
rect 895 192 908 194
rect 859 189 861 192
rect 869 189 871 192
rect 879 189 881 192
rect 895 189 897 192
rect 822 182 828 183
rect 822 178 823 182
rect 827 178 828 182
rect 822 177 828 178
rect 869 167 871 171
rect 879 167 881 171
rect 811 158 813 162
rect 859 158 861 162
rect 906 183 908 192
rect 961 190 963 201
rect 969 196 971 210
rect 981 199 983 207
rect 977 198 983 199
rect 969 193 973 196
rect 977 194 978 198
rect 982 194 983 198
rect 977 193 983 194
rect 971 190 973 193
rect 981 190 983 193
rect 906 182 912 183
rect 906 178 907 182
rect 911 178 912 182
rect 906 177 912 178
rect 961 175 963 180
rect 971 175 973 180
rect 967 174 973 175
rect 967 170 968 174
rect 972 170 973 174
rect 981 173 983 178
rect 967 169 973 170
rect 895 158 897 162
rect 128 148 130 152
rect 52 140 58 141
rect 42 132 44 137
rect 52 136 53 140
rect 57 136 58 140
rect 52 135 58 136
rect 52 130 54 135
rect 62 130 64 135
rect 113 132 119 133
rect 113 128 114 132
rect 118 128 119 132
rect 113 127 119 128
rect 42 117 44 120
rect 52 117 54 120
rect 42 116 48 117
rect 42 112 43 116
rect 47 112 48 116
rect 52 114 56 117
rect 42 111 48 112
rect 42 103 44 111
rect 54 100 56 114
rect 62 109 64 120
rect 117 118 119 127
rect 164 148 166 152
rect 212 148 214 152
rect 144 139 146 143
rect 154 139 156 143
rect 197 132 203 133
rect 197 128 198 132
rect 202 128 203 132
rect 197 127 203 128
rect 128 118 130 121
rect 144 118 146 121
rect 154 118 156 121
rect 164 118 166 121
rect 117 116 130 118
rect 136 116 146 118
rect 150 117 156 118
rect 61 108 67 109
rect 120 108 122 116
rect 136 112 138 116
rect 150 113 151 117
rect 155 113 156 117
rect 150 112 156 113
rect 160 117 166 118
rect 160 113 161 117
rect 165 113 166 117
rect 201 118 203 127
rect 248 148 250 152
rect 228 139 230 143
rect 238 139 240 143
rect 284 140 290 141
rect 274 132 276 137
rect 284 136 285 140
rect 289 136 290 140
rect 484 140 486 144
rect 284 135 290 136
rect 212 118 214 121
rect 228 118 230 121
rect 238 118 240 121
rect 248 118 250 121
rect 284 130 286 135
rect 294 130 296 135
rect 408 132 414 133
rect 398 124 400 129
rect 408 128 409 132
rect 413 128 414 132
rect 408 127 414 128
rect 201 116 214 118
rect 220 116 230 118
rect 234 117 240 118
rect 160 112 166 113
rect 129 111 138 112
rect 61 104 62 108
rect 66 104 67 108
rect 61 103 67 104
rect 61 100 63 103
rect 42 93 44 97
rect 129 107 130 111
rect 134 107 138 111
rect 154 108 156 112
rect 129 106 138 107
rect 136 103 138 106
rect 146 103 148 108
rect 154 106 158 108
rect 156 103 158 106
rect 163 103 165 112
rect 204 108 206 116
rect 220 112 222 116
rect 234 113 235 117
rect 239 113 240 117
rect 234 112 240 113
rect 244 117 250 118
rect 244 113 245 117
rect 249 113 250 117
rect 244 112 250 113
rect 274 117 276 120
rect 284 117 286 120
rect 274 116 280 117
rect 274 112 275 116
rect 279 112 280 116
rect 284 114 288 117
rect 213 111 222 112
rect 120 96 122 99
rect 120 94 125 96
rect 54 86 56 91
rect 61 86 63 91
rect 123 86 125 94
rect 136 90 138 94
rect 146 86 148 94
rect 213 107 214 111
rect 218 107 222 111
rect 238 108 240 112
rect 213 106 222 107
rect 220 103 222 106
rect 230 103 232 108
rect 238 106 242 108
rect 240 103 242 106
rect 247 103 249 112
rect 274 111 280 112
rect 274 103 276 111
rect 204 96 206 99
rect 204 94 209 96
rect 156 86 158 91
rect 163 86 165 91
rect 123 84 148 86
rect 207 86 209 94
rect 220 90 222 94
rect 230 86 232 94
rect 286 100 288 114
rect 294 109 296 120
rect 408 122 410 127
rect 418 122 420 127
rect 469 124 475 125
rect 469 120 470 124
rect 474 120 475 124
rect 469 119 475 120
rect 398 109 400 112
rect 408 109 410 112
rect 293 108 299 109
rect 293 104 294 108
rect 298 104 299 108
rect 293 103 299 104
rect 398 108 404 109
rect 398 104 399 108
rect 403 104 404 108
rect 408 106 412 109
rect 398 103 404 104
rect 293 100 295 103
rect 274 93 276 97
rect 398 95 400 103
rect 240 86 242 91
rect 247 86 249 91
rect 207 84 232 86
rect 286 86 288 91
rect 293 86 295 91
rect 410 92 412 106
rect 418 101 420 112
rect 473 110 475 119
rect 520 140 522 144
rect 568 140 570 144
rect 500 131 502 135
rect 510 131 512 135
rect 553 124 559 125
rect 553 120 554 124
rect 558 120 559 124
rect 553 119 559 120
rect 484 110 486 113
rect 500 110 502 113
rect 510 110 512 113
rect 520 110 522 113
rect 473 108 486 110
rect 492 108 502 110
rect 506 109 512 110
rect 417 100 423 101
rect 476 100 478 108
rect 492 104 494 108
rect 506 105 507 109
rect 511 105 512 109
rect 506 104 512 105
rect 516 109 522 110
rect 516 105 517 109
rect 521 105 522 109
rect 557 110 559 119
rect 604 140 606 144
rect 584 131 586 135
rect 594 131 596 135
rect 844 142 846 146
rect 768 134 774 135
rect 640 132 646 133
rect 630 124 632 129
rect 640 128 641 132
rect 645 128 646 132
rect 640 127 646 128
rect 568 110 570 113
rect 584 110 586 113
rect 594 110 596 113
rect 604 110 606 113
rect 640 122 642 127
rect 650 122 652 127
rect 758 126 760 131
rect 768 130 769 134
rect 773 130 774 134
rect 768 129 774 130
rect 768 124 770 129
rect 778 124 780 129
rect 829 126 835 127
rect 829 122 830 126
rect 834 122 835 126
rect 829 121 835 122
rect 557 108 570 110
rect 576 108 586 110
rect 590 109 596 110
rect 516 104 522 105
rect 485 103 494 104
rect 417 96 418 100
rect 422 96 423 100
rect 417 95 423 96
rect 417 92 419 95
rect 398 85 400 89
rect 485 99 486 103
rect 490 99 494 103
rect 510 100 512 104
rect 485 98 494 99
rect 492 95 494 98
rect 502 95 504 100
rect 510 98 514 100
rect 512 95 514 98
rect 519 95 521 104
rect 560 100 562 108
rect 576 104 578 108
rect 590 105 591 109
rect 595 105 596 109
rect 590 104 596 105
rect 600 109 606 110
rect 600 105 601 109
rect 605 105 606 109
rect 600 104 606 105
rect 630 109 632 112
rect 640 109 642 112
rect 630 108 636 109
rect 630 104 631 108
rect 635 104 636 108
rect 640 106 644 109
rect 569 103 578 104
rect 476 88 478 91
rect 476 86 481 88
rect 39 79 41 83
rect 50 79 52 83
rect 57 79 59 83
rect 39 56 41 65
rect 77 73 79 78
rect 87 73 89 78
rect 97 76 99 81
rect 107 79 109 83
rect 410 78 412 83
rect 417 78 419 83
rect 479 78 481 86
rect 492 82 494 86
rect 502 78 504 86
rect 569 99 570 103
rect 574 99 578 103
rect 594 100 596 104
rect 569 98 578 99
rect 576 95 578 98
rect 586 95 588 100
rect 594 98 598 100
rect 596 95 598 98
rect 603 95 605 104
rect 630 103 636 104
rect 630 95 632 103
rect 560 88 562 91
rect 560 86 565 88
rect 512 78 514 83
rect 519 78 521 83
rect 479 76 504 78
rect 563 78 565 86
rect 576 82 578 86
rect 586 78 588 86
rect 642 92 644 106
rect 650 101 652 112
rect 758 111 760 114
rect 768 111 770 114
rect 758 110 764 111
rect 758 106 759 110
rect 763 106 764 110
rect 768 108 772 111
rect 758 105 764 106
rect 649 100 655 101
rect 649 96 650 100
rect 654 96 655 100
rect 758 97 760 105
rect 649 95 655 96
rect 649 92 651 95
rect 630 85 632 89
rect 770 94 772 108
rect 778 103 780 114
rect 833 112 835 121
rect 880 142 882 146
rect 928 142 930 146
rect 860 133 862 137
rect 870 133 872 137
rect 913 126 919 127
rect 913 122 914 126
rect 918 122 919 126
rect 913 121 919 122
rect 844 112 846 115
rect 860 112 862 115
rect 870 112 872 115
rect 880 112 882 115
rect 833 110 846 112
rect 852 110 862 112
rect 866 111 872 112
rect 777 102 783 103
rect 836 102 838 110
rect 852 106 854 110
rect 866 107 867 111
rect 871 107 872 111
rect 866 106 872 107
rect 876 111 882 112
rect 876 107 877 111
rect 881 107 882 111
rect 917 112 919 121
rect 964 142 966 146
rect 944 133 946 137
rect 954 133 956 137
rect 1000 134 1006 135
rect 990 126 992 131
rect 1000 130 1001 134
rect 1005 130 1006 134
rect 1000 129 1006 130
rect 928 112 930 115
rect 944 112 946 115
rect 954 112 956 115
rect 964 112 966 115
rect 1000 124 1002 129
rect 1010 124 1012 129
rect 917 110 930 112
rect 936 110 946 112
rect 950 111 956 112
rect 876 106 882 107
rect 845 105 854 106
rect 777 98 778 102
rect 782 98 783 102
rect 777 97 783 98
rect 777 94 779 97
rect 758 87 760 91
rect 845 101 846 105
rect 850 101 854 105
rect 870 102 872 106
rect 845 100 854 101
rect 852 97 854 100
rect 862 97 864 102
rect 870 100 874 102
rect 872 97 874 100
rect 879 97 881 106
rect 920 102 922 110
rect 936 106 938 110
rect 950 107 951 111
rect 955 107 956 111
rect 950 106 956 107
rect 960 111 966 112
rect 960 107 961 111
rect 965 107 966 111
rect 960 106 966 107
rect 990 111 992 114
rect 1000 111 1002 114
rect 990 110 996 111
rect 990 106 991 110
rect 995 106 996 110
rect 1000 108 1004 111
rect 929 105 938 106
rect 836 90 838 93
rect 836 88 841 90
rect 596 78 598 83
rect 603 78 605 83
rect 563 76 588 78
rect 642 78 644 83
rect 649 78 651 83
rect 770 80 772 85
rect 777 80 779 85
rect 839 80 841 88
rect 852 84 854 88
rect 862 80 864 88
rect 929 101 930 105
rect 934 101 938 105
rect 954 102 956 106
rect 929 100 938 101
rect 936 97 938 100
rect 946 97 948 102
rect 954 100 958 102
rect 956 97 958 100
rect 963 97 965 106
rect 990 105 996 106
rect 990 97 992 105
rect 920 90 922 93
rect 920 88 925 90
rect 872 80 874 85
rect 879 80 881 85
rect 839 78 864 80
rect 923 80 925 88
rect 936 84 938 88
rect 946 80 948 88
rect 1002 94 1004 108
rect 1010 103 1012 114
rect 1009 102 1015 103
rect 1009 98 1010 102
rect 1014 98 1015 102
rect 1009 97 1015 98
rect 1009 94 1011 97
rect 990 87 992 91
rect 956 80 958 85
rect 963 80 965 85
rect 923 78 948 80
rect 1002 80 1004 85
rect 1009 80 1011 85
rect 135 69 137 73
rect 145 69 147 73
rect 155 69 157 73
rect 50 56 52 59
rect 57 56 59 59
rect 77 56 79 59
rect 87 56 89 59
rect 37 55 43 56
rect 37 51 38 55
rect 42 51 43 55
rect 37 50 43 51
rect 47 55 53 56
rect 47 51 48 55
rect 52 51 53 55
rect 47 50 53 51
rect 57 55 79 56
rect 57 51 58 55
rect 62 51 65 55
rect 69 51 79 55
rect 57 50 79 51
rect 83 55 89 56
rect 83 51 84 55
rect 88 51 89 55
rect 83 50 89 51
rect 97 53 99 66
rect 107 63 109 66
rect 103 62 109 63
rect 103 58 104 62
rect 108 58 109 62
rect 103 57 109 58
rect 97 52 103 53
rect 39 47 41 50
rect 49 47 51 50
rect 59 47 61 50
rect 72 47 74 50
rect 77 47 79 50
rect 84 47 86 50
rect 97 49 98 52
rect 94 48 98 49
rect 102 48 103 52
rect 94 47 103 48
rect 94 44 96 47
rect 107 44 109 57
rect 135 55 137 63
rect 131 54 137 55
rect 145 54 147 63
rect 155 54 157 63
rect 491 61 493 65
rect 501 61 503 65
rect 511 61 513 65
rect 851 63 853 67
rect 861 63 863 67
rect 871 63 873 67
rect 131 50 132 54
rect 136 50 137 54
rect 151 53 157 54
rect 131 49 137 50
rect 94 26 96 31
rect 135 36 137 49
rect 145 47 147 50
rect 151 49 152 53
rect 156 49 157 53
rect 151 48 157 49
rect 141 46 147 47
rect 141 42 142 46
rect 146 42 147 46
rect 141 41 147 42
rect 142 36 144 41
rect 155 39 157 48
rect 491 47 493 55
rect 487 46 493 47
rect 501 46 503 55
rect 511 46 513 55
rect 851 49 853 57
rect 487 42 488 46
rect 492 42 493 46
rect 507 45 513 46
rect 487 41 493 42
rect 39 17 41 19
rect 49 17 51 19
rect 59 1 61 19
rect 72 17 74 19
rect 77 17 79 19
rect 84 -1 86 19
rect 107 15 109 19
rect 491 28 493 41
rect 501 39 503 42
rect 507 41 508 45
rect 512 41 513 45
rect 847 48 853 49
rect 861 48 863 57
rect 871 48 873 57
rect 847 44 848 48
rect 852 44 853 48
rect 867 47 873 48
rect 847 43 853 44
rect 507 40 513 41
rect 497 38 503 39
rect 497 34 498 38
rect 502 34 503 38
rect 497 33 503 34
rect 498 28 500 33
rect 511 31 513 40
rect 155 23 157 27
rect 135 14 137 18
rect 142 14 144 18
rect 851 30 853 43
rect 861 41 863 44
rect 867 43 868 47
rect 872 43 873 47
rect 867 42 873 43
rect 857 40 863 41
rect 857 36 858 40
rect 862 36 863 40
rect 857 35 863 36
rect 858 30 860 35
rect 871 33 873 42
rect 511 15 513 19
rect 871 17 873 21
rect 491 6 493 10
rect 498 6 500 10
rect 851 8 853 12
rect 858 8 860 12
<< ndiffusion >>
rect 750 245 755 252
rect 501 244 508 245
rect 501 240 502 244
rect 506 240 508 244
rect 501 239 508 240
rect 510 244 518 245
rect 510 240 512 244
rect 516 240 518 244
rect 510 239 518 240
rect 520 244 528 245
rect 520 240 522 244
rect 526 240 528 244
rect 520 239 528 240
rect 530 244 537 245
rect 530 240 532 244
rect 536 240 537 244
rect 530 239 537 240
rect 728 244 735 245
rect 728 240 729 244
rect 733 240 735 244
rect 728 239 735 240
rect 730 232 735 239
rect 737 240 745 245
rect 737 236 739 240
rect 743 236 745 240
rect 737 235 745 236
rect 747 243 755 245
rect 747 239 749 243
rect 753 239 755 243
rect 747 238 755 239
rect 757 251 765 252
rect 757 247 759 251
rect 763 247 765 251
rect 757 238 765 247
rect 767 251 774 252
rect 767 247 769 251
rect 773 247 774 251
rect 767 244 774 247
rect 780 245 785 252
rect 767 240 769 244
rect 773 240 774 244
rect 767 238 774 240
rect 778 244 785 245
rect 778 240 779 244
rect 783 240 785 244
rect 778 239 785 240
rect 747 235 752 238
rect 737 232 742 235
rect 780 232 785 239
rect 787 232 792 252
rect 794 246 801 252
rect 861 246 868 247
rect 794 237 803 246
rect 794 233 796 237
rect 800 233 803 237
rect 794 232 803 233
rect 805 244 812 246
rect 805 240 807 244
rect 811 240 812 244
rect 861 242 862 246
rect 866 242 868 246
rect 861 241 868 242
rect 870 246 878 247
rect 870 242 872 246
rect 876 242 878 246
rect 870 241 878 242
rect 880 246 888 247
rect 880 242 882 246
rect 886 242 888 246
rect 880 241 888 242
rect 890 246 897 247
rect 890 242 892 246
rect 896 242 897 246
rect 890 241 897 242
rect 805 239 812 240
rect 805 232 810 239
rect 741 224 747 225
rect 381 222 387 223
rect 381 218 382 222
rect 386 218 387 222
rect 381 217 387 218
rect 408 222 414 223
rect 408 218 409 222
rect 413 218 414 222
rect 408 217 414 218
rect 365 214 370 217
rect 363 213 370 214
rect 363 209 364 213
rect 368 209 370 213
rect 363 208 370 209
rect 372 208 377 217
rect 379 211 387 217
rect 379 208 389 211
rect 381 205 389 208
rect 391 210 398 211
rect 391 206 393 210
rect 397 206 398 210
rect 391 205 398 206
rect 408 205 416 217
rect 418 205 423 217
rect 425 214 430 217
rect 492 222 498 223
rect 492 218 493 222
rect 497 218 498 222
rect 492 217 498 218
rect 425 212 433 214
rect 425 208 427 212
rect 431 208 433 212
rect 425 205 433 208
rect 435 210 443 214
rect 435 206 437 210
rect 441 206 443 210
rect 435 205 443 206
rect 445 213 454 214
rect 445 209 449 213
rect 453 209 454 213
rect 445 205 459 209
rect 454 200 459 205
rect 461 206 466 209
rect 461 205 468 206
rect 492 205 500 217
rect 502 205 507 217
rect 509 214 514 217
rect 613 222 619 223
rect 613 218 614 222
rect 618 218 619 222
rect 613 217 619 218
rect 741 220 742 224
rect 746 220 747 224
rect 741 219 747 220
rect 768 224 774 225
rect 768 220 769 224
rect 773 220 774 224
rect 768 219 774 220
rect 597 214 602 217
rect 509 212 517 214
rect 509 208 511 212
rect 515 208 517 212
rect 509 205 517 208
rect 519 210 527 214
rect 519 206 521 210
rect 525 206 527 210
rect 519 205 527 206
rect 529 213 538 214
rect 529 209 533 213
rect 537 209 538 213
rect 595 213 602 214
rect 595 209 596 213
rect 600 209 602 213
rect 529 205 543 209
rect 461 201 463 205
rect 467 201 468 205
rect 461 200 468 201
rect 538 200 543 205
rect 545 206 550 209
rect 595 208 602 209
rect 604 208 609 217
rect 611 211 619 217
rect 725 216 730 219
rect 723 215 730 216
rect 723 211 724 215
rect 728 211 730 215
rect 611 208 621 211
rect 545 205 552 206
rect 545 201 547 205
rect 551 201 552 205
rect 545 200 552 201
rect 613 205 621 208
rect 623 210 630 211
rect 723 210 730 211
rect 732 210 737 219
rect 739 213 747 219
rect 739 210 749 213
rect 623 206 625 210
rect 629 206 630 210
rect 623 205 630 206
rect 741 207 749 210
rect 751 212 758 213
rect 751 208 753 212
rect 757 208 758 212
rect 751 207 758 208
rect 768 207 776 219
rect 778 207 783 219
rect 785 216 790 219
rect 852 224 858 225
rect 852 220 853 224
rect 857 220 858 224
rect 852 219 858 220
rect 785 214 793 216
rect 785 210 787 214
rect 791 210 793 214
rect 785 207 793 210
rect 795 212 803 216
rect 795 208 797 212
rect 801 208 803 212
rect 795 207 803 208
rect 805 215 814 216
rect 805 211 809 215
rect 813 211 814 215
rect 805 207 819 211
rect 814 202 819 207
rect 821 208 826 211
rect 821 207 828 208
rect 852 207 860 219
rect 862 207 867 219
rect 869 216 874 219
rect 973 224 979 225
rect 973 220 974 224
rect 978 220 979 224
rect 973 219 979 220
rect 957 216 962 219
rect 869 214 877 216
rect 869 210 871 214
rect 875 210 877 214
rect 869 207 877 210
rect 879 212 887 216
rect 879 208 881 212
rect 885 208 887 212
rect 879 207 887 208
rect 889 215 898 216
rect 889 211 893 215
rect 897 211 898 215
rect 955 215 962 216
rect 955 211 956 215
rect 960 211 962 215
rect 889 207 903 211
rect 821 203 823 207
rect 827 203 828 207
rect 821 202 828 203
rect 898 202 903 207
rect 905 208 910 211
rect 955 210 962 211
rect 964 210 969 219
rect 971 213 979 219
rect 971 210 981 213
rect 905 207 912 208
rect 905 203 907 207
rect 911 203 912 207
rect 905 202 912 203
rect 973 207 981 210
rect 983 212 990 213
rect 983 208 985 212
rect 989 208 990 212
rect 983 207 990 208
rect 35 102 42 103
rect 35 98 36 102
rect 40 98 42 102
rect 35 97 42 98
rect 44 100 52 103
rect 113 107 120 108
rect 113 103 114 107
rect 118 103 120 107
rect 113 102 120 103
rect 44 97 54 100
rect 46 91 54 97
rect 56 91 61 100
rect 63 99 70 100
rect 115 99 120 102
rect 122 103 127 108
rect 197 107 204 108
rect 197 103 198 107
rect 202 103 204 107
rect 122 99 136 103
rect 63 95 65 99
rect 69 95 70 99
rect 63 94 70 95
rect 127 95 128 99
rect 132 95 136 99
rect 127 94 136 95
rect 138 102 146 103
rect 138 98 140 102
rect 144 98 146 102
rect 138 94 146 98
rect 148 100 156 103
rect 148 96 150 100
rect 154 96 156 100
rect 148 94 156 96
rect 63 91 68 94
rect 46 90 52 91
rect 46 86 47 90
rect 51 86 52 90
rect 46 85 52 86
rect 151 91 156 94
rect 158 91 163 103
rect 165 91 173 103
rect 197 102 204 103
rect 199 99 204 102
rect 206 103 211 108
rect 206 99 220 103
rect 211 95 212 99
rect 216 95 220 99
rect 211 94 220 95
rect 222 102 230 103
rect 222 98 224 102
rect 228 98 230 102
rect 222 94 230 98
rect 232 100 240 103
rect 232 96 234 100
rect 238 96 240 100
rect 232 94 240 96
rect 167 90 173 91
rect 167 86 168 90
rect 172 86 173 90
rect 167 85 173 86
rect 235 91 240 94
rect 242 91 247 103
rect 249 91 257 103
rect 267 102 274 103
rect 267 98 268 102
rect 272 98 274 102
rect 267 97 274 98
rect 276 100 284 103
rect 276 97 286 100
rect 278 91 286 97
rect 288 91 293 100
rect 295 99 302 100
rect 295 95 297 99
rect 301 95 302 99
rect 295 94 302 95
rect 391 94 398 95
rect 295 91 300 94
rect 251 90 257 91
rect 251 86 252 90
rect 256 86 257 90
rect 251 85 257 86
rect 278 90 284 91
rect 278 86 279 90
rect 283 86 284 90
rect 391 90 392 94
rect 396 90 398 94
rect 391 89 398 90
rect 400 92 408 95
rect 469 99 476 100
rect 469 95 470 99
rect 474 95 476 99
rect 469 94 476 95
rect 400 89 410 92
rect 278 85 284 86
rect 402 83 410 89
rect 412 83 417 92
rect 419 91 426 92
rect 471 91 476 94
rect 478 95 483 100
rect 553 99 560 100
rect 553 95 554 99
rect 558 95 560 99
rect 478 91 492 95
rect 419 87 421 91
rect 425 87 426 91
rect 419 86 426 87
rect 483 87 484 91
rect 488 87 492 91
rect 483 86 492 87
rect 494 94 502 95
rect 494 90 496 94
rect 500 90 502 94
rect 494 86 502 90
rect 504 92 512 95
rect 504 88 506 92
rect 510 88 512 92
rect 504 86 512 88
rect 419 83 424 86
rect 34 72 39 79
rect 32 71 39 72
rect 32 67 33 71
rect 37 67 39 71
rect 32 65 39 67
rect 41 78 50 79
rect 41 74 44 78
rect 48 74 50 78
rect 41 65 50 74
rect 43 59 50 65
rect 52 59 57 79
rect 59 72 64 79
rect 102 76 107 79
rect 92 73 97 76
rect 59 71 66 72
rect 59 67 61 71
rect 65 67 66 71
rect 59 66 66 67
rect 70 71 77 73
rect 70 67 71 71
rect 75 67 77 71
rect 59 59 64 66
rect 70 64 77 67
rect 70 60 71 64
rect 75 60 77 64
rect 70 59 77 60
rect 79 64 87 73
rect 79 60 81 64
rect 85 60 87 64
rect 79 59 87 60
rect 89 72 97 73
rect 89 68 91 72
rect 95 68 97 72
rect 89 66 97 68
rect 99 75 107 76
rect 99 71 101 75
rect 105 71 107 75
rect 99 66 107 71
rect 109 72 114 79
rect 402 82 408 83
rect 402 78 403 82
rect 407 78 408 82
rect 402 77 408 78
rect 507 83 512 86
rect 514 83 519 95
rect 521 83 529 95
rect 553 94 560 95
rect 555 91 560 94
rect 562 95 567 100
rect 562 91 576 95
rect 567 87 568 91
rect 572 87 576 91
rect 567 86 576 87
rect 578 94 586 95
rect 578 90 580 94
rect 584 90 586 94
rect 578 86 586 90
rect 588 92 596 95
rect 588 88 590 92
rect 594 88 596 92
rect 588 86 596 88
rect 523 82 529 83
rect 523 78 524 82
rect 528 78 529 82
rect 523 77 529 78
rect 591 83 596 86
rect 598 83 603 95
rect 605 83 613 95
rect 623 94 630 95
rect 623 90 624 94
rect 628 90 630 94
rect 623 89 630 90
rect 632 92 640 95
rect 751 96 758 97
rect 751 92 752 96
rect 756 92 758 96
rect 632 89 642 92
rect 634 83 642 89
rect 644 83 649 92
rect 651 91 658 92
rect 751 91 758 92
rect 760 94 768 97
rect 829 101 836 102
rect 829 97 830 101
rect 834 97 836 101
rect 829 96 836 97
rect 760 91 770 94
rect 651 87 653 91
rect 657 87 658 91
rect 651 86 658 87
rect 651 83 656 86
rect 762 85 770 91
rect 772 85 777 94
rect 779 93 786 94
rect 831 93 836 96
rect 838 97 843 102
rect 913 101 920 102
rect 913 97 914 101
rect 918 97 920 101
rect 838 93 852 97
rect 779 89 781 93
rect 785 89 786 93
rect 779 88 786 89
rect 843 89 844 93
rect 848 89 852 93
rect 843 88 852 89
rect 854 96 862 97
rect 854 92 856 96
rect 860 92 862 96
rect 854 88 862 92
rect 864 94 872 97
rect 864 90 866 94
rect 870 90 872 94
rect 864 88 872 90
rect 779 85 784 88
rect 607 82 613 83
rect 607 78 608 82
rect 612 78 613 82
rect 607 77 613 78
rect 634 82 640 83
rect 634 78 635 82
rect 639 78 640 82
rect 762 84 768 85
rect 762 80 763 84
rect 767 80 768 84
rect 762 79 768 80
rect 867 85 872 88
rect 874 85 879 97
rect 881 85 889 97
rect 913 96 920 97
rect 915 93 920 96
rect 922 97 927 102
rect 922 93 936 97
rect 927 89 928 93
rect 932 89 936 93
rect 927 88 936 89
rect 938 96 946 97
rect 938 92 940 96
rect 944 92 946 96
rect 938 88 946 92
rect 948 94 956 97
rect 948 90 950 94
rect 954 90 956 94
rect 948 88 956 90
rect 883 84 889 85
rect 883 80 884 84
rect 888 80 889 84
rect 883 79 889 80
rect 951 85 956 88
rect 958 85 963 97
rect 965 85 973 97
rect 983 96 990 97
rect 983 92 984 96
rect 988 92 990 96
rect 983 91 990 92
rect 992 94 1000 97
rect 992 91 1002 94
rect 994 85 1002 91
rect 1004 85 1009 94
rect 1011 93 1018 94
rect 1011 89 1013 93
rect 1017 89 1018 93
rect 1011 88 1018 89
rect 1011 85 1016 88
rect 967 84 973 85
rect 967 80 968 84
rect 972 80 973 84
rect 967 79 973 80
rect 994 84 1000 85
rect 994 80 995 84
rect 999 80 1000 84
rect 994 79 1000 80
rect 634 77 640 78
rect 109 71 116 72
rect 109 67 111 71
rect 115 67 116 71
rect 109 66 116 67
rect 128 68 135 69
rect 89 59 94 66
rect 128 64 129 68
rect 133 64 135 68
rect 128 63 135 64
rect 137 68 145 69
rect 137 64 139 68
rect 143 64 145 68
rect 137 63 145 64
rect 147 68 155 69
rect 147 64 149 68
rect 153 64 155 68
rect 147 63 155 64
rect 157 68 164 69
rect 157 64 159 68
rect 163 64 164 68
rect 157 63 164 64
rect 844 62 851 63
rect 484 60 491 61
rect 484 56 485 60
rect 489 56 491 60
rect 484 55 491 56
rect 493 60 501 61
rect 493 56 495 60
rect 499 56 501 60
rect 493 55 501 56
rect 503 60 511 61
rect 503 56 505 60
rect 509 56 511 60
rect 503 55 511 56
rect 513 60 520 61
rect 513 56 515 60
rect 519 56 520 60
rect 844 58 845 62
rect 849 58 851 62
rect 844 57 851 58
rect 853 62 861 63
rect 853 58 855 62
rect 859 58 861 62
rect 853 57 861 58
rect 863 62 871 63
rect 863 58 865 62
rect 869 58 871 62
rect 863 57 871 58
rect 873 62 880 63
rect 873 58 875 62
rect 879 58 880 62
rect 873 57 880 58
rect 513 55 520 56
<< pdiffusion >>
rect 512 289 521 290
rect 512 285 514 289
rect 518 285 521 289
rect 512 281 521 285
rect 501 280 508 281
rect 501 276 502 280
rect 506 276 508 280
rect 501 275 508 276
rect 503 269 508 275
rect 510 272 521 281
rect 523 272 528 290
rect 530 283 535 290
rect 530 282 537 283
rect 530 278 532 282
rect 536 278 537 282
rect 730 280 735 292
rect 530 277 537 278
rect 728 279 735 280
rect 530 272 535 277
rect 728 275 729 279
rect 733 275 735 279
rect 728 272 735 275
rect 510 269 518 272
rect 728 268 729 272
rect 733 268 735 272
rect 728 267 735 268
rect 737 291 746 292
rect 737 287 740 291
rect 744 287 746 291
rect 769 291 783 292
rect 769 289 775 291
rect 737 280 746 287
rect 753 280 758 289
rect 737 267 748 280
rect 750 272 758 280
rect 750 268 752 272
rect 756 268 758 272
rect 750 267 758 268
rect 753 264 758 267
rect 760 264 765 289
rect 767 287 775 289
rect 779 287 783 291
rect 767 284 783 287
rect 767 280 775 284
rect 779 280 783 284
rect 767 264 783 280
rect 785 283 793 292
rect 785 279 787 283
rect 791 279 793 283
rect 785 276 793 279
rect 785 272 787 276
rect 791 272 793 276
rect 785 264 793 272
rect 795 291 803 292
rect 795 287 797 291
rect 801 287 803 291
rect 795 284 803 287
rect 795 280 797 284
rect 801 280 803 284
rect 795 264 803 280
rect 805 277 810 292
rect 872 291 881 292
rect 872 287 874 291
rect 878 287 881 291
rect 872 283 881 287
rect 861 282 868 283
rect 861 278 862 282
rect 866 278 868 282
rect 861 277 868 278
rect 805 276 812 277
rect 805 272 807 276
rect 811 272 812 276
rect 805 269 812 272
rect 863 271 868 277
rect 870 274 881 283
rect 883 274 888 292
rect 890 285 895 292
rect 890 284 897 285
rect 890 280 892 284
rect 896 280 897 284
rect 890 279 897 280
rect 890 274 895 279
rect 870 271 878 274
rect 805 265 807 269
rect 811 265 812 269
rect 805 264 812 265
rect 362 183 369 188
rect 362 179 363 183
rect 367 179 369 183
rect 362 178 369 179
rect 371 187 379 188
rect 371 183 373 187
rect 377 183 379 187
rect 371 178 379 183
rect 381 187 389 188
rect 381 183 383 187
rect 387 183 389 187
rect 381 178 389 183
rect 383 176 389 178
rect 391 187 398 188
rect 391 183 393 187
rect 397 183 398 187
rect 391 182 398 183
rect 391 176 396 182
rect 410 172 415 187
rect 408 171 415 172
rect 408 167 409 171
rect 413 167 415 171
rect 408 166 415 167
rect 410 160 415 166
rect 417 179 425 187
rect 417 175 419 179
rect 423 175 425 179
rect 417 169 425 175
rect 427 186 435 187
rect 427 182 429 186
rect 433 182 435 186
rect 427 169 435 182
rect 437 172 451 187
rect 437 169 445 172
rect 417 160 422 169
rect 439 168 445 169
rect 449 168 451 172
rect 439 165 451 168
rect 439 161 445 165
rect 449 161 451 165
rect 439 160 451 161
rect 453 186 460 187
rect 453 182 455 186
rect 459 182 460 186
rect 453 181 460 182
rect 453 160 458 181
rect 494 172 499 187
rect 492 171 499 172
rect 492 167 493 171
rect 497 167 499 171
rect 492 166 499 167
rect 494 160 499 166
rect 501 179 509 187
rect 501 175 503 179
rect 507 175 509 179
rect 501 169 509 175
rect 511 186 519 187
rect 511 182 513 186
rect 517 182 519 186
rect 511 169 519 182
rect 521 172 535 187
rect 521 169 529 172
rect 501 160 506 169
rect 523 168 529 169
rect 533 168 535 172
rect 523 165 535 168
rect 523 161 529 165
rect 533 161 535 165
rect 523 160 535 161
rect 537 186 544 187
rect 537 182 539 186
rect 543 182 544 186
rect 537 181 544 182
rect 594 183 601 188
rect 537 160 542 181
rect 594 179 595 183
rect 599 179 601 183
rect 594 178 601 179
rect 603 187 611 188
rect 603 183 605 187
rect 609 183 611 187
rect 603 178 611 183
rect 613 187 621 188
rect 613 183 615 187
rect 619 183 621 187
rect 613 178 621 183
rect 615 176 621 178
rect 623 187 630 188
rect 623 183 625 187
rect 629 183 630 187
rect 623 182 630 183
rect 722 185 729 190
rect 623 176 628 182
rect 722 181 723 185
rect 727 181 729 185
rect 722 180 729 181
rect 731 189 739 190
rect 731 185 733 189
rect 737 185 739 189
rect 731 180 739 185
rect 741 189 749 190
rect 741 185 743 189
rect 747 185 749 189
rect 741 180 749 185
rect 743 178 749 180
rect 751 189 758 190
rect 751 185 753 189
rect 757 185 758 189
rect 751 184 758 185
rect 751 178 756 184
rect 770 174 775 189
rect 768 173 775 174
rect 768 169 769 173
rect 773 169 775 173
rect 768 168 775 169
rect 770 162 775 168
rect 777 181 785 189
rect 777 177 779 181
rect 783 177 785 181
rect 777 171 785 177
rect 787 188 795 189
rect 787 184 789 188
rect 793 184 795 188
rect 787 171 795 184
rect 797 174 811 189
rect 797 171 805 174
rect 777 162 782 171
rect 799 170 805 171
rect 809 170 811 174
rect 799 167 811 170
rect 799 163 805 167
rect 809 163 811 167
rect 799 162 811 163
rect 813 188 820 189
rect 813 184 815 188
rect 819 184 820 188
rect 813 183 820 184
rect 813 162 818 183
rect 854 174 859 189
rect 852 173 859 174
rect 852 169 853 173
rect 857 169 859 173
rect 852 168 859 169
rect 854 162 859 168
rect 861 181 869 189
rect 861 177 863 181
rect 867 177 869 181
rect 861 171 869 177
rect 871 188 879 189
rect 871 184 873 188
rect 877 184 879 188
rect 871 171 879 184
rect 881 174 895 189
rect 881 171 889 174
rect 861 162 866 171
rect 883 170 889 171
rect 893 170 895 174
rect 883 167 895 170
rect 883 163 889 167
rect 893 163 895 167
rect 883 162 895 163
rect 897 188 904 189
rect 897 184 899 188
rect 903 184 904 188
rect 897 183 904 184
rect 954 185 961 190
rect 897 162 902 183
rect 954 181 955 185
rect 959 181 961 185
rect 954 180 961 181
rect 963 189 971 190
rect 963 185 965 189
rect 969 185 971 189
rect 963 180 971 185
rect 973 189 981 190
rect 973 185 975 189
rect 979 185 981 189
rect 973 180 981 185
rect 975 178 981 180
rect 983 189 990 190
rect 983 185 985 189
rect 989 185 990 189
rect 983 184 990 185
rect 983 178 988 184
rect 37 126 42 132
rect 35 125 42 126
rect 35 121 36 125
rect 40 121 42 125
rect 35 120 42 121
rect 44 130 50 132
rect 44 125 52 130
rect 44 121 46 125
rect 50 121 52 125
rect 44 120 52 121
rect 54 125 62 130
rect 54 121 56 125
rect 60 121 62 125
rect 54 120 62 121
rect 64 129 71 130
rect 64 125 66 129
rect 70 125 71 129
rect 123 127 128 148
rect 64 120 71 125
rect 121 126 128 127
rect 121 122 122 126
rect 126 122 128 126
rect 121 121 128 122
rect 130 147 142 148
rect 130 143 132 147
rect 136 143 142 147
rect 130 140 142 143
rect 130 136 132 140
rect 136 139 142 140
rect 159 139 164 148
rect 136 136 144 139
rect 130 121 144 136
rect 146 126 154 139
rect 146 122 148 126
rect 152 122 154 126
rect 146 121 154 122
rect 156 133 164 139
rect 156 129 158 133
rect 162 129 164 133
rect 156 121 164 129
rect 166 142 171 148
rect 166 141 173 142
rect 166 137 168 141
rect 172 137 173 141
rect 166 136 173 137
rect 166 121 171 136
rect 207 127 212 148
rect 205 126 212 127
rect 205 122 206 126
rect 210 122 212 126
rect 205 121 212 122
rect 214 147 226 148
rect 214 143 216 147
rect 220 143 226 147
rect 214 140 226 143
rect 214 136 216 140
rect 220 139 226 140
rect 243 139 248 148
rect 220 136 228 139
rect 214 121 228 136
rect 230 126 238 139
rect 230 122 232 126
rect 236 122 238 126
rect 230 121 238 122
rect 240 133 248 139
rect 240 129 242 133
rect 246 129 248 133
rect 240 121 248 129
rect 250 142 255 148
rect 250 141 257 142
rect 250 137 252 141
rect 256 137 257 141
rect 250 136 257 137
rect 250 121 255 136
rect 269 126 274 132
rect 267 125 274 126
rect 267 121 268 125
rect 272 121 274 125
rect 267 120 274 121
rect 276 130 282 132
rect 276 125 284 130
rect 276 121 278 125
rect 282 121 284 125
rect 276 120 284 121
rect 286 125 294 130
rect 286 121 288 125
rect 292 121 294 125
rect 286 120 294 121
rect 296 129 303 130
rect 296 125 298 129
rect 302 125 303 129
rect 296 120 303 125
rect 393 118 398 124
rect 391 117 398 118
rect 391 113 392 117
rect 396 113 398 117
rect 391 112 398 113
rect 400 122 406 124
rect 400 117 408 122
rect 400 113 402 117
rect 406 113 408 117
rect 400 112 408 113
rect 410 117 418 122
rect 410 113 412 117
rect 416 113 418 117
rect 410 112 418 113
rect 420 121 427 122
rect 420 117 422 121
rect 426 117 427 121
rect 479 119 484 140
rect 420 112 427 117
rect 477 118 484 119
rect 477 114 478 118
rect 482 114 484 118
rect 477 113 484 114
rect 486 139 498 140
rect 486 135 488 139
rect 492 135 498 139
rect 486 132 498 135
rect 486 128 488 132
rect 492 131 498 132
rect 515 131 520 140
rect 492 128 500 131
rect 486 113 500 128
rect 502 118 510 131
rect 502 114 504 118
rect 508 114 510 118
rect 502 113 510 114
rect 512 125 520 131
rect 512 121 514 125
rect 518 121 520 125
rect 512 113 520 121
rect 522 134 527 140
rect 522 133 529 134
rect 522 129 524 133
rect 528 129 529 133
rect 522 128 529 129
rect 522 113 527 128
rect 563 119 568 140
rect 561 118 568 119
rect 561 114 562 118
rect 566 114 568 118
rect 561 113 568 114
rect 570 139 582 140
rect 570 135 572 139
rect 576 135 582 139
rect 570 132 582 135
rect 570 128 572 132
rect 576 131 582 132
rect 599 131 604 140
rect 576 128 584 131
rect 570 113 584 128
rect 586 118 594 131
rect 586 114 588 118
rect 592 114 594 118
rect 586 113 594 114
rect 596 125 604 131
rect 596 121 598 125
rect 602 121 604 125
rect 596 113 604 121
rect 606 134 611 140
rect 606 133 613 134
rect 606 129 608 133
rect 612 129 613 133
rect 606 128 613 129
rect 606 113 611 128
rect 625 118 630 124
rect 623 117 630 118
rect 623 113 624 117
rect 628 113 630 117
rect 623 112 630 113
rect 632 122 638 124
rect 632 117 640 122
rect 632 113 634 117
rect 638 113 640 117
rect 632 112 640 113
rect 642 117 650 122
rect 642 113 644 117
rect 648 113 650 117
rect 642 112 650 113
rect 652 121 659 122
rect 652 117 654 121
rect 658 117 659 121
rect 753 120 758 126
rect 652 112 659 117
rect 751 119 758 120
rect 751 115 752 119
rect 756 115 758 119
rect 751 114 758 115
rect 760 124 766 126
rect 760 119 768 124
rect 760 115 762 119
rect 766 115 768 119
rect 760 114 768 115
rect 770 119 778 124
rect 770 115 772 119
rect 776 115 778 119
rect 770 114 778 115
rect 780 123 787 124
rect 780 119 782 123
rect 786 119 787 123
rect 839 121 844 142
rect 780 114 787 119
rect 837 120 844 121
rect 837 116 838 120
rect 842 116 844 120
rect 837 115 844 116
rect 846 141 858 142
rect 846 137 848 141
rect 852 137 858 141
rect 846 134 858 137
rect 846 130 848 134
rect 852 133 858 134
rect 875 133 880 142
rect 852 130 860 133
rect 846 115 860 130
rect 862 120 870 133
rect 862 116 864 120
rect 868 116 870 120
rect 862 115 870 116
rect 872 127 880 133
rect 872 123 874 127
rect 878 123 880 127
rect 872 115 880 123
rect 882 136 887 142
rect 882 135 889 136
rect 882 131 884 135
rect 888 131 889 135
rect 882 130 889 131
rect 882 115 887 130
rect 923 121 928 142
rect 921 120 928 121
rect 921 116 922 120
rect 926 116 928 120
rect 921 115 928 116
rect 930 141 942 142
rect 930 137 932 141
rect 936 137 942 141
rect 930 134 942 137
rect 930 130 932 134
rect 936 133 942 134
rect 959 133 964 142
rect 936 130 944 133
rect 930 115 944 130
rect 946 120 954 133
rect 946 116 948 120
rect 952 116 954 120
rect 946 115 954 116
rect 956 127 964 133
rect 956 123 958 127
rect 962 123 964 127
rect 956 115 964 123
rect 966 136 971 142
rect 966 135 973 136
rect 966 131 968 135
rect 972 131 973 135
rect 966 130 973 131
rect 966 115 971 130
rect 985 120 990 126
rect 983 119 990 120
rect 983 115 984 119
rect 988 115 990 119
rect 983 114 990 115
rect 992 124 998 126
rect 992 119 1000 124
rect 992 115 994 119
rect 998 115 1000 119
rect 992 114 1000 115
rect 1002 119 1010 124
rect 1002 115 1004 119
rect 1008 115 1010 119
rect 1002 114 1010 115
rect 1012 123 1019 124
rect 1012 119 1014 123
rect 1018 119 1019 123
rect 1012 114 1019 119
rect 32 46 39 47
rect 32 42 33 46
rect 37 42 39 46
rect 32 39 39 42
rect 32 35 33 39
rect 37 35 39 39
rect 32 34 39 35
rect 34 19 39 34
rect 41 31 49 47
rect 41 27 43 31
rect 47 27 49 31
rect 41 24 49 27
rect 41 20 43 24
rect 47 20 49 24
rect 41 19 49 20
rect 51 39 59 47
rect 51 35 53 39
rect 57 35 59 39
rect 51 32 59 35
rect 51 28 53 32
rect 57 28 59 32
rect 51 19 59 28
rect 61 31 72 47
rect 61 27 65 31
rect 69 27 72 31
rect 61 24 72 27
rect 61 20 65 24
rect 69 20 72 24
rect 61 19 72 20
rect 74 19 77 47
rect 79 19 84 47
rect 86 44 91 47
rect 86 43 94 44
rect 86 39 88 43
rect 92 39 94 43
rect 86 31 94 39
rect 96 31 107 44
rect 86 19 91 31
rect 98 24 107 31
rect 98 20 100 24
rect 104 20 107 24
rect 98 19 107 20
rect 109 43 116 44
rect 109 39 111 43
rect 115 39 116 43
rect 109 36 116 39
rect 147 36 155 39
rect 109 32 111 36
rect 115 32 116 36
rect 109 31 116 32
rect 130 31 135 36
rect 109 19 114 31
rect 128 30 135 31
rect 128 26 129 30
rect 133 26 135 30
rect 128 25 135 26
rect 130 18 135 25
rect 137 18 142 36
rect 144 27 155 36
rect 157 33 162 39
rect 157 32 164 33
rect 157 28 159 32
rect 163 28 164 32
rect 503 28 511 31
rect 157 27 164 28
rect 144 23 153 27
rect 486 23 491 28
rect 144 19 147 23
rect 151 19 153 23
rect 484 22 491 23
rect 144 18 153 19
rect 484 18 485 22
rect 489 18 491 22
rect 484 17 491 18
rect 486 10 491 17
rect 493 10 498 28
rect 500 19 511 28
rect 513 25 518 31
rect 863 30 871 33
rect 846 25 851 30
rect 513 24 520 25
rect 513 20 515 24
rect 519 20 520 24
rect 513 19 520 20
rect 844 24 851 25
rect 844 20 845 24
rect 849 20 851 24
rect 844 19 851 20
rect 500 15 509 19
rect 500 11 503 15
rect 507 11 509 15
rect 500 10 509 11
rect 846 12 851 19
rect 853 12 858 30
rect 860 21 871 30
rect 873 27 878 33
rect 873 26 880 27
rect 873 22 875 26
rect 879 22 880 26
rect 873 21 880 22
rect 860 17 869 21
rect 860 13 863 17
rect 867 13 869 17
rect 860 12 869 13
<< metal1 >>
rect 261 381 264 382
rect 261 378 1054 381
rect 261 254 264 378
rect 339 361 1061 364
rect 339 290 342 361
rect 685 345 1061 348
rect 682 301 685 344
rect 758 313 761 324
rect 850 311 853 328
rect 901 298 1025 299
rect 724 297 824 298
rect 857 297 1025 298
rect 541 296 670 297
rect 497 294 670 296
rect 691 295 1025 297
rect 691 294 901 295
rect 497 293 863 294
rect 497 292 541 293
rect 497 288 503 292
rect 507 289 541 292
rect 507 288 514 289
rect 513 285 514 288
rect 518 288 541 289
rect 660 291 863 293
rect 518 285 519 288
rect 501 280 514 282
rect 501 276 502 280
rect 506 278 514 280
rect 517 278 532 282
rect 536 278 537 282
rect 501 275 506 276
rect 501 258 505 275
rect 517 274 521 278
rect 501 245 505 254
rect 509 270 521 274
rect 525 272 542 275
rect 509 259 513 270
rect 525 266 529 272
rect 660 273 665 291
rect 724 290 740 291
rect 739 287 740 290
rect 744 290 775 291
rect 744 287 745 290
rect 774 287 775 290
rect 779 290 797 291
rect 779 287 780 290
rect 774 284 780 287
rect 796 287 797 290
rect 801 290 824 291
rect 857 290 863 291
rect 867 291 901 294
rect 867 290 874 291
rect 801 287 802 290
rect 873 287 874 290
rect 878 290 901 291
rect 878 287 879 290
rect 796 284 802 287
rect 728 280 741 284
rect 774 280 775 284
rect 779 280 780 284
rect 787 283 791 284
rect 728 279 733 280
rect 728 275 729 279
rect 744 276 768 280
rect 796 280 797 284
rect 801 280 802 284
rect 861 282 874 284
rect 787 276 791 279
rect 807 276 813 277
rect 516 262 519 266
rect 523 262 529 266
rect 509 251 513 255
rect 524 254 529 258
rect 533 253 537 263
rect 624 254 646 257
rect 509 247 526 251
rect -4 241 429 244
rect 501 244 506 245
rect 522 244 526 247
rect 501 240 502 244
rect 501 237 506 240
rect 511 240 512 244
rect 516 240 517 244
rect -4 232 430 235
rect 511 232 517 240
rect 522 239 526 240
rect 531 240 532 244
rect 536 240 537 244
rect 531 232 537 240
rect 497 228 503 232
rect 507 228 531 232
rect 535 228 541 232
rect 497 226 541 228
rect 358 224 631 226
rect 324 222 631 224
rect 324 219 382 222
rect 261 161 264 210
rect 1 153 313 154
rect 1 151 311 153
rect 1 150 256 151
rect 1 146 37 150
rect 41 146 51 150
rect 55 146 65 150
rect 69 147 148 150
rect 69 146 132 147
rect 1 35 5 146
rect 35 126 39 133
rect 35 125 40 126
rect 35 121 36 125
rect 43 125 47 146
rect 50 140 63 141
rect 50 136 53 140
rect 57 136 59 140
rect 50 135 63 136
rect 50 128 56 135
rect 66 129 70 146
rect 136 146 148 147
rect 152 147 232 150
rect 152 146 216 147
rect 113 135 125 141
rect 132 140 136 143
rect 220 146 232 147
rect 236 146 256 150
rect 267 150 311 151
rect 146 137 168 141
rect 172 137 173 141
rect 197 140 209 141
rect 182 137 202 140
rect 146 136 150 137
rect 132 135 136 136
rect 113 132 118 135
rect 43 121 46 125
rect 50 121 51 125
rect 55 121 56 125
rect 60 121 61 125
rect 66 124 70 125
rect 113 131 114 132
rect 109 128 114 131
rect 139 132 150 136
rect 139 128 143 132
rect 157 129 158 133
rect 162 129 173 133
rect 35 120 40 121
rect 35 112 39 120
rect 55 116 61 121
rect 42 112 43 116
rect 47 112 61 116
rect 67 114 71 117
rect 105 114 108 128
rect 113 127 118 128
rect 122 126 143 128
rect 35 103 39 108
rect 35 102 40 103
rect 35 98 36 102
rect 40 98 47 101
rect 35 95 47 98
rect 51 99 55 112
rect 114 122 122 123
rect 126 124 143 126
rect 114 119 126 122
rect 67 108 71 110
rect 58 104 62 108
rect 66 104 71 108
rect 58 103 71 104
rect 114 107 118 119
rect 139 117 143 124
rect 147 122 148 126
rect 152 125 153 126
rect 152 122 164 125
rect 147 121 164 122
rect 160 118 164 121
rect 160 117 165 118
rect 128 111 134 116
rect 139 113 151 117
rect 155 113 156 117
rect 160 113 161 117
rect 128 109 130 111
rect 121 107 130 109
rect 160 112 165 113
rect 169 113 173 129
rect 160 108 164 112
rect 121 103 134 107
rect 140 104 164 108
rect 169 109 171 113
rect 114 102 118 103
rect 140 102 144 104
rect 51 95 65 99
rect 69 95 70 99
rect 127 95 128 99
rect 132 95 133 99
rect 169 100 173 109
rect 140 97 144 98
rect 149 96 150 100
rect 154 96 173 100
rect 182 97 185 137
rect 197 136 202 137
rect 206 136 209 140
rect 197 135 209 136
rect 216 140 220 143
rect 267 146 269 150
rect 273 146 283 150
rect 287 146 297 150
rect 301 148 311 150
rect 301 146 307 148
rect 230 137 252 141
rect 256 137 257 141
rect 230 136 234 137
rect 216 135 220 136
rect 197 132 202 135
rect 197 128 198 132
rect 223 132 234 136
rect 223 128 227 132
rect 241 129 242 133
rect 246 129 257 133
rect 197 127 202 128
rect 206 126 227 128
rect 198 122 206 123
rect 210 124 227 126
rect 198 119 210 122
rect 198 107 202 119
rect 223 117 227 124
rect 231 122 232 126
rect 236 125 237 126
rect 236 122 248 125
rect 231 121 248 122
rect 244 118 248 121
rect 253 121 257 129
rect 260 121 263 144
rect 253 118 263 121
rect 267 126 271 133
rect 267 125 272 126
rect 267 121 268 125
rect 275 125 279 146
rect 282 140 295 141
rect 282 136 285 140
rect 289 136 291 140
rect 282 135 295 136
rect 282 128 288 135
rect 298 129 302 146
rect 275 121 278 125
rect 282 121 283 125
rect 287 121 288 125
rect 292 121 293 125
rect 298 124 302 125
rect 267 120 272 121
rect 244 117 249 118
rect 212 111 218 116
rect 223 113 235 117
rect 239 113 240 117
rect 244 113 245 117
rect 212 109 214 111
rect 205 107 214 109
rect 244 112 249 113
rect 244 108 248 112
rect 205 103 218 107
rect 224 104 248 108
rect 198 102 202 103
rect 224 102 228 104
rect 127 90 133 95
rect 211 95 212 99
rect 216 95 217 99
rect 253 100 257 118
rect 267 112 271 120
rect 287 116 293 121
rect 274 112 275 116
rect 279 112 293 116
rect 299 115 303 117
rect 224 97 228 98
rect 233 96 234 100
rect 238 96 257 100
rect 261 109 271 112
rect 261 97 264 109
rect 211 90 217 95
rect 267 103 271 109
rect 267 102 272 103
rect 267 98 268 102
rect 272 98 279 101
rect 267 95 279 98
rect 283 99 287 112
rect 299 108 303 111
rect 290 104 294 108
rect 298 104 303 108
rect 290 103 303 104
rect 324 103 330 219
rect 358 218 382 219
rect 386 218 392 222
rect 396 218 409 222
rect 413 218 462 222
rect 466 218 493 222
rect 497 218 546 222
rect 550 218 614 222
rect 618 218 624 222
rect 628 218 631 222
rect 363 209 364 213
rect 368 209 382 213
rect 362 204 375 205
rect 362 200 367 204
rect 371 200 375 204
rect 362 197 366 200
rect 378 196 382 209
rect 386 210 398 213
rect 386 207 393 210
rect 397 206 398 210
rect 393 205 398 206
rect 394 199 398 205
rect 448 213 454 218
rect 401 199 404 211
rect 394 196 404 199
rect 408 208 427 212
rect 431 208 432 212
rect 437 210 441 211
rect 362 191 366 193
rect 372 192 386 196
rect 390 192 391 196
rect 372 187 378 192
rect 394 188 398 196
rect 393 187 398 188
rect 363 183 367 184
rect 372 183 373 187
rect 377 183 378 187
rect 382 183 383 187
rect 387 183 390 187
rect 363 162 367 179
rect 377 173 383 180
rect 370 172 383 173
rect 374 168 376 172
rect 380 168 383 172
rect 370 167 383 168
rect 386 162 390 183
rect 397 183 398 187
rect 393 182 398 183
rect 394 175 398 182
rect 408 179 412 208
rect 448 209 449 213
rect 453 209 454 213
rect 532 213 538 218
rect 492 208 511 212
rect 515 208 516 212
rect 521 210 525 211
rect 437 204 441 206
rect 463 205 467 206
rect 417 200 441 204
rect 447 201 460 205
rect 417 196 421 200
rect 416 195 421 196
rect 451 199 460 201
rect 451 197 453 199
rect 420 191 421 195
rect 425 191 426 195
rect 430 191 442 195
rect 447 192 453 197
rect 416 190 421 191
rect 417 187 421 190
rect 417 186 434 187
rect 417 183 429 186
rect 428 182 429 183
rect 433 182 434 186
rect 438 184 442 191
rect 463 189 467 201
rect 492 199 496 208
rect 532 209 533 213
rect 537 209 538 213
rect 595 209 596 213
rect 600 209 614 213
rect 521 204 525 206
rect 547 205 551 206
rect 494 195 496 199
rect 501 200 525 204
rect 531 201 544 205
rect 501 196 505 200
rect 455 186 467 189
rect 438 182 455 184
rect 459 185 467 186
rect 438 180 459 182
rect 463 180 468 181
rect 408 175 419 179
rect 423 175 424 179
rect 438 176 442 180
rect 431 172 442 176
rect 467 176 468 180
rect 463 173 468 176
rect 492 179 496 195
rect 500 195 505 196
rect 535 199 544 201
rect 535 197 537 199
rect 504 191 505 195
rect 509 191 510 195
rect 514 191 526 195
rect 531 192 537 197
rect 500 190 505 191
rect 501 187 505 190
rect 501 186 518 187
rect 501 183 513 186
rect 512 182 513 183
rect 517 182 518 186
rect 522 184 526 191
rect 547 189 551 201
rect 594 204 607 205
rect 594 200 599 204
rect 603 200 607 204
rect 594 198 598 200
rect 539 186 551 189
rect 522 182 539 184
rect 543 185 551 186
rect 610 196 614 209
rect 618 210 630 213
rect 618 207 625 210
rect 629 206 630 210
rect 625 205 630 206
rect 626 200 630 205
rect 522 180 543 182
rect 547 180 552 181
rect 557 180 560 194
rect 594 191 598 194
rect 604 192 618 196
rect 622 192 623 196
rect 604 187 610 192
rect 626 188 630 196
rect 625 187 630 188
rect 492 175 503 179
rect 507 175 508 179
rect 522 176 526 180
rect 445 172 449 173
rect 431 171 435 172
rect 408 167 409 171
rect 413 167 435 171
rect 445 165 449 168
rect 456 172 468 173
rect 456 168 459 172
rect 463 168 468 172
rect 515 172 526 176
rect 551 177 560 180
rect 595 183 599 184
rect 604 183 605 187
rect 609 183 610 187
rect 614 183 615 187
rect 619 183 622 187
rect 551 176 552 177
rect 547 173 552 176
rect 529 172 533 173
rect 515 171 519 172
rect 456 167 468 168
rect 492 167 493 171
rect 497 167 519 171
rect 358 158 364 162
rect 368 158 378 162
rect 382 158 392 162
rect 396 158 429 162
rect 433 161 445 162
rect 529 165 533 168
rect 540 167 552 173
rect 449 161 513 162
rect 433 158 513 161
rect 517 161 529 162
rect 595 162 599 179
rect 609 173 615 180
rect 602 172 615 173
rect 606 168 608 172
rect 612 168 615 172
rect 602 167 615 168
rect 618 162 622 183
rect 629 183 630 187
rect 625 182 630 183
rect 626 175 630 182
rect 660 162 664 273
rect 728 272 733 275
rect 728 268 729 272
rect 728 267 733 268
rect 742 272 748 276
rect 752 272 756 273
rect 764 272 787 276
rect 791 272 804 276
rect 728 245 732 267
rect 742 263 746 272
rect 742 258 746 259
rect 749 264 756 268
rect 759 264 797 268
rect 749 253 753 264
rect 759 261 764 264
rect 756 260 764 261
rect 792 260 796 264
rect 760 256 764 260
rect 772 256 775 260
rect 779 256 782 260
rect 786 256 789 260
rect 756 255 764 256
rect 735 249 736 253
rect 740 251 753 253
rect 769 251 773 252
rect 740 249 759 251
rect 749 247 759 249
rect 763 247 764 251
rect 776 247 780 256
rect 792 255 796 256
rect 800 261 804 272
rect 811 272 813 276
rect 807 269 813 272
rect 811 265 813 269
rect 807 264 813 265
rect 800 260 806 261
rect 800 256 802 260
rect 800 255 806 256
rect 800 252 804 255
rect 784 248 804 252
rect 728 244 733 245
rect 728 240 729 244
rect 769 244 773 247
rect 784 244 788 248
rect 809 244 813 264
rect 728 239 733 240
rect 739 240 743 241
rect 748 239 749 243
rect 753 240 769 243
rect 778 240 779 244
rect 783 240 788 244
rect 791 240 807 244
rect 811 240 813 244
rect 753 239 773 240
rect 739 234 743 236
rect 795 234 796 237
rect 724 233 796 234
rect 800 234 801 237
rect 838 236 841 280
rect 861 278 862 282
rect 866 280 874 282
rect 877 280 892 284
rect 896 280 897 284
rect 861 277 866 278
rect 861 247 865 277
rect 877 276 881 280
rect 869 272 881 276
rect 885 274 902 277
rect 869 261 873 272
rect 885 268 889 274
rect 876 264 879 268
rect 883 264 889 268
rect 869 253 873 257
rect 884 256 889 260
rect 893 255 897 265
rect 928 260 931 286
rect 1020 275 1025 295
rect 869 249 886 253
rect 922 249 1001 252
rect 861 246 866 247
rect 882 246 886 249
rect 861 242 862 246
rect 861 239 866 242
rect 871 242 872 246
rect 876 242 877 246
rect 800 233 824 234
rect 724 228 824 233
rect 871 234 877 242
rect 882 241 886 242
rect 891 242 892 246
rect 896 242 897 246
rect 891 234 897 242
rect 904 240 1001 243
rect 1005 240 1007 243
rect 857 230 863 234
rect 867 230 891 234
rect 895 230 901 234
rect 857 228 901 230
rect 718 226 991 228
rect 533 161 596 162
rect 517 158 596 161
rect 600 158 610 162
rect 614 158 624 162
rect 628 158 664 162
rect 358 154 664 158
rect 358 148 359 154
rect 365 148 664 154
rect 358 146 664 148
rect 357 144 664 146
rect 684 224 991 226
rect 684 221 742 224
rect 357 142 663 144
rect 357 138 393 142
rect 397 138 407 142
rect 411 138 421 142
rect 425 139 504 142
rect 425 138 488 139
rect 283 95 297 99
rect 301 95 302 99
rect 329 98 330 103
rect 34 86 37 90
rect 41 86 47 90
rect 51 86 115 90
rect 119 86 168 90
rect 172 86 199 90
rect 203 86 252 90
rect 256 86 269 90
rect 273 86 279 90
rect 283 86 307 90
rect 34 85 307 86
rect 20 82 307 85
rect 20 78 120 82
rect 20 77 44 78
rect 43 74 44 77
rect 48 77 120 78
rect 124 80 168 82
rect 48 74 49 77
rect 101 75 105 77
rect 124 76 130 80
rect 134 76 158 80
rect 162 76 168 80
rect 71 71 91 72
rect 0 15 5 35
rect 31 67 33 71
rect 37 67 44 71
rect 48 67 53 71
rect 56 67 61 71
rect 65 67 66 71
rect 75 68 91 71
rect 95 68 96 72
rect 101 70 105 71
rect 111 71 116 72
rect 31 47 35 67
rect 56 63 60 67
rect 71 64 75 67
rect 115 67 116 71
rect 111 66 116 67
rect 40 59 60 63
rect 40 56 44 59
rect 38 55 44 56
rect 42 51 44 55
rect 38 50 44 51
rect 31 46 37 47
rect 31 42 33 46
rect 31 39 37 42
rect 31 35 33 39
rect 40 39 44 50
rect 48 55 52 56
rect 64 55 68 64
rect 80 60 81 64
rect 85 62 95 64
rect 85 60 104 62
rect 71 59 75 60
rect 91 58 104 60
rect 108 58 109 62
rect 80 55 88 56
rect 55 51 58 55
rect 62 51 65 55
rect 69 51 70 55
rect 80 51 84 55
rect 48 47 52 51
rect 80 50 88 51
rect 80 47 85 50
rect 91 47 95 58
rect 47 43 85 47
rect 88 43 95 47
rect 98 52 102 53
rect 98 39 102 48
rect 112 44 116 66
rect 128 68 134 76
rect 128 64 129 68
rect 133 64 134 68
rect 139 68 143 69
rect 148 68 154 76
rect 148 64 149 68
rect 153 64 154 68
rect 159 68 164 71
rect 163 64 164 68
rect 139 61 143 64
rect 159 63 164 64
rect 139 57 156 61
rect 40 35 53 39
rect 57 35 80 39
rect 88 38 92 39
rect 96 35 102 39
rect 111 43 116 44
rect 115 39 116 43
rect 128 45 132 55
rect 136 50 141 54
rect 152 53 156 57
rect 136 42 142 46
rect 146 42 149 46
rect 111 36 116 39
rect 31 34 37 35
rect 53 32 57 35
rect 42 27 43 31
rect 47 27 48 31
rect 76 31 100 35
rect 115 32 116 36
rect 136 36 140 42
rect 152 38 156 49
rect 123 33 140 36
rect 144 34 156 38
rect 160 58 164 63
rect 160 52 279 58
rect 111 31 116 32
rect 53 27 57 28
rect 64 27 65 31
rect 69 27 70 31
rect 103 30 116 31
rect 144 30 148 34
rect 160 33 164 52
rect 276 46 279 52
rect 159 32 164 33
rect 103 29 117 30
rect 103 27 115 29
rect 42 24 48 27
rect 42 21 43 24
rect 20 20 43 21
rect 47 21 48 24
rect 64 24 70 27
rect 114 25 115 27
rect 119 25 121 28
rect 128 26 129 30
rect 133 26 148 30
rect 151 28 159 30
rect 163 28 164 32
rect 151 26 164 28
rect 301 29 306 82
rect 345 80 350 123
rect 301 24 343 29
rect 348 24 349 29
rect 357 27 361 138
rect 391 118 395 125
rect 391 117 396 118
rect 391 113 392 117
rect 399 117 403 138
rect 406 132 419 133
rect 406 128 409 132
rect 413 128 415 132
rect 406 127 419 128
rect 406 120 412 127
rect 422 121 426 138
rect 492 138 504 139
rect 508 139 588 142
rect 508 138 572 139
rect 469 127 481 133
rect 488 132 492 135
rect 576 138 588 139
rect 592 138 625 142
rect 629 138 639 142
rect 643 138 653 142
rect 657 138 663 142
rect 502 129 524 133
rect 528 129 529 133
rect 502 128 506 129
rect 488 127 492 128
rect 469 124 474 127
rect 469 123 470 124
rect 461 120 470 123
rect 495 124 506 128
rect 495 120 499 124
rect 513 121 514 125
rect 518 121 529 125
rect 399 113 402 117
rect 406 113 407 117
rect 411 113 412 117
rect 416 113 417 117
rect 422 116 426 117
rect 391 112 396 113
rect 391 104 395 112
rect 411 108 417 113
rect 398 104 399 108
rect 403 104 417 108
rect 423 106 427 109
rect 391 95 395 100
rect 391 94 396 95
rect 391 90 392 94
rect 396 90 403 93
rect 391 87 403 90
rect 407 91 411 104
rect 423 100 427 102
rect 414 96 418 100
rect 422 96 427 100
rect 414 95 427 96
rect 451 98 455 112
rect 461 106 464 120
rect 469 119 474 120
rect 478 118 499 120
rect 470 114 478 115
rect 482 116 499 118
rect 470 111 482 114
rect 470 99 474 111
rect 495 109 499 116
rect 503 114 504 118
rect 508 117 509 118
rect 508 114 520 117
rect 503 113 520 114
rect 516 110 520 113
rect 516 109 521 110
rect 484 103 490 108
rect 495 105 507 109
rect 511 105 512 109
rect 516 105 517 109
rect 484 101 486 103
rect 477 99 486 101
rect 516 104 521 105
rect 525 105 529 121
rect 516 100 520 104
rect 477 95 490 99
rect 496 96 520 100
rect 525 101 527 105
rect 470 94 474 95
rect 496 94 500 96
rect 407 87 421 91
rect 425 87 426 91
rect 483 87 484 91
rect 488 87 489 91
rect 525 92 529 101
rect 496 89 500 90
rect 505 88 506 92
rect 510 88 529 92
rect 539 90 542 129
rect 553 132 565 133
rect 553 128 558 132
rect 562 128 565 132
rect 553 127 565 128
rect 572 132 576 135
rect 586 129 608 133
rect 612 129 613 133
rect 586 128 590 129
rect 572 127 576 128
rect 553 124 558 127
rect 553 120 554 124
rect 579 124 590 128
rect 579 120 583 124
rect 597 121 598 125
rect 602 121 613 125
rect 553 119 558 120
rect 562 118 583 120
rect 554 114 562 115
rect 566 116 583 118
rect 554 111 566 114
rect 554 99 558 111
rect 579 109 583 116
rect 587 114 588 118
rect 592 117 593 118
rect 592 114 604 117
rect 587 113 604 114
rect 600 110 604 113
rect 609 114 613 121
rect 623 118 627 125
rect 623 117 628 118
rect 609 111 616 114
rect 623 113 624 117
rect 631 117 635 138
rect 638 132 651 133
rect 638 128 641 132
rect 645 128 647 132
rect 638 127 651 128
rect 638 120 644 127
rect 654 121 658 138
rect 631 113 634 117
rect 638 113 639 117
rect 643 113 644 117
rect 648 113 649 117
rect 654 116 658 117
rect 623 112 628 113
rect 600 109 605 110
rect 568 103 574 108
rect 579 105 591 109
rect 595 105 596 109
rect 600 105 601 109
rect 568 101 570 103
rect 561 99 570 101
rect 600 104 605 105
rect 600 100 604 104
rect 561 95 574 99
rect 580 96 604 100
rect 554 94 558 95
rect 580 94 584 96
rect 483 82 489 87
rect 567 87 568 91
rect 572 87 573 91
rect 609 92 613 111
rect 623 104 627 112
rect 643 108 649 113
rect 630 104 631 108
rect 635 104 649 108
rect 655 107 659 109
rect 580 89 584 90
rect 589 88 590 92
rect 594 88 613 92
rect 617 101 627 104
rect 617 89 620 101
rect 539 85 542 86
rect 567 82 573 87
rect 623 95 627 101
rect 623 94 628 95
rect 623 90 624 94
rect 628 90 635 93
rect 623 87 635 90
rect 639 91 643 104
rect 684 105 690 221
rect 718 220 742 221
rect 746 220 752 224
rect 756 220 769 224
rect 773 220 822 224
rect 826 220 853 224
rect 857 220 906 224
rect 910 220 974 224
rect 978 220 984 224
rect 988 220 991 224
rect 723 211 724 215
rect 728 211 742 215
rect 722 206 735 207
rect 722 202 727 206
rect 731 202 735 206
rect 722 199 726 202
rect 738 198 742 211
rect 746 212 758 215
rect 746 209 753 212
rect 757 208 758 212
rect 753 207 758 208
rect 754 201 758 207
rect 808 215 814 220
rect 761 201 764 213
rect 754 198 764 201
rect 768 210 787 214
rect 791 210 792 214
rect 797 212 801 213
rect 722 193 726 195
rect 732 194 746 198
rect 750 194 751 198
rect 732 189 738 194
rect 754 190 758 198
rect 753 189 758 190
rect 768 189 772 210
rect 808 211 809 215
rect 813 211 814 215
rect 836 213 841 217
rect 892 215 898 220
rect 797 206 801 208
rect 823 207 827 208
rect 777 202 801 206
rect 807 203 820 207
rect 777 198 781 202
rect 776 197 781 198
rect 811 201 820 203
rect 811 199 813 201
rect 780 193 781 197
rect 785 193 786 197
rect 790 193 802 197
rect 807 194 813 199
rect 776 192 781 193
rect 723 185 727 186
rect 732 185 733 189
rect 737 185 738 189
rect 742 185 743 189
rect 747 185 750 189
rect 723 164 727 181
rect 737 175 743 182
rect 730 174 743 175
rect 734 170 736 174
rect 740 170 743 174
rect 730 169 743 170
rect 746 164 750 185
rect 757 185 758 189
rect 766 185 772 189
rect 777 189 781 192
rect 777 188 794 189
rect 777 185 789 188
rect 753 184 758 185
rect 754 177 758 184
rect 768 181 772 185
rect 788 184 789 185
rect 793 184 794 188
rect 798 186 802 193
rect 823 191 827 203
rect 815 188 827 191
rect 838 190 841 213
rect 852 210 871 214
rect 875 210 876 214
rect 881 212 885 213
rect 852 201 856 210
rect 892 211 893 215
rect 897 211 898 215
rect 955 211 956 215
rect 960 211 974 215
rect 881 206 885 208
rect 907 207 911 208
rect 854 197 856 201
rect 861 202 885 206
rect 891 203 904 207
rect 861 198 865 202
rect 798 184 815 186
rect 819 187 827 188
rect 798 182 819 184
rect 823 182 828 183
rect 768 177 779 181
rect 783 177 784 181
rect 798 178 802 182
rect 791 174 802 178
rect 827 178 828 182
rect 823 175 828 178
rect 852 181 856 197
rect 860 197 865 198
rect 895 201 904 203
rect 895 199 897 201
rect 864 193 865 197
rect 869 193 870 197
rect 874 193 886 197
rect 891 194 897 199
rect 860 192 865 193
rect 861 189 865 192
rect 861 188 878 189
rect 861 185 873 188
rect 872 184 873 185
rect 877 184 878 188
rect 882 186 886 193
rect 907 191 911 203
rect 954 206 967 207
rect 954 202 959 206
rect 963 202 967 206
rect 954 200 958 202
rect 899 188 911 191
rect 882 184 899 186
rect 903 187 911 188
rect 970 198 974 211
rect 978 212 990 215
rect 978 209 985 212
rect 989 208 990 212
rect 985 207 990 208
rect 986 202 990 207
rect 882 182 903 184
rect 907 182 912 183
rect 917 182 920 196
rect 954 193 958 196
rect 964 194 978 198
rect 982 194 983 198
rect 964 189 970 194
rect 986 190 990 198
rect 985 189 990 190
rect 852 177 863 181
rect 867 177 868 181
rect 882 178 886 182
rect 805 174 809 175
rect 791 173 795 174
rect 768 169 769 173
rect 773 169 795 173
rect 805 167 809 170
rect 816 174 828 175
rect 816 170 819 174
rect 823 170 828 174
rect 875 174 886 178
rect 911 179 920 182
rect 955 185 959 186
rect 964 185 965 189
rect 969 185 970 189
rect 974 185 975 189
rect 979 185 982 189
rect 911 178 912 179
rect 907 175 912 178
rect 889 174 893 175
rect 875 173 879 174
rect 816 169 828 170
rect 852 169 853 173
rect 857 169 879 173
rect 718 160 724 164
rect 728 160 738 164
rect 742 160 752 164
rect 756 160 789 164
rect 793 163 805 164
rect 889 167 893 170
rect 900 169 912 175
rect 809 163 873 164
rect 793 160 873 163
rect 877 163 889 164
rect 955 164 959 181
rect 969 175 975 182
rect 962 174 975 175
rect 966 170 968 174
rect 972 170 975 174
rect 962 169 975 170
rect 978 164 982 185
rect 989 185 990 189
rect 985 184 990 185
rect 986 177 990 184
rect 1020 164 1024 275
rect 893 163 956 164
rect 877 160 956 163
rect 960 160 970 164
rect 974 160 984 164
rect 988 160 1024 164
rect 718 148 1024 160
rect 655 100 659 103
rect 646 96 650 100
rect 654 96 659 100
rect 646 95 659 96
rect 682 98 683 103
rect 689 100 690 105
rect 717 146 1024 148
rect 717 144 1023 146
rect 717 140 753 144
rect 757 140 767 144
rect 771 140 781 144
rect 785 141 864 144
rect 785 140 848 141
rect 639 87 653 91
rect 657 87 658 91
rect 390 78 393 82
rect 397 78 403 82
rect 407 78 471 82
rect 475 78 524 82
rect 528 78 555 82
rect 559 78 608 82
rect 612 78 625 82
rect 629 78 635 82
rect 639 80 663 82
rect 682 80 688 98
rect 639 78 693 80
rect 373 76 693 78
rect 376 75 693 76
rect 376 74 663 75
rect 376 68 454 74
rect 480 72 524 74
rect 480 68 486 72
rect 490 68 514 72
rect 518 68 524 72
rect 393 28 398 68
rect 484 60 490 68
rect 484 56 485 60
rect 489 56 490 60
rect 495 60 499 61
rect 504 60 510 68
rect 504 56 505 60
rect 509 56 510 60
rect 515 60 520 63
rect 519 56 520 60
rect 495 53 499 56
rect 515 55 520 56
rect 495 49 512 53
rect 64 21 65 24
rect 47 20 65 21
rect 69 21 70 24
rect 99 21 100 24
rect 69 20 100 21
rect 104 21 105 24
rect 104 20 120 21
rect 146 20 147 23
rect 20 18 120 20
rect 18 15 120 18
rect 124 19 147 20
rect 151 20 152 23
rect 151 19 158 20
rect 124 16 158 19
rect 162 16 168 20
rect 124 15 168 16
rect 0 12 168 15
rect 0 11 124 12
rect 356 7 361 27
rect 452 26 455 47
rect 484 37 488 47
rect 492 42 497 46
rect 508 45 512 49
rect 492 34 498 38
rect 502 34 505 38
rect 492 28 496 34
rect 508 30 512 41
rect 479 25 496 28
rect 500 26 512 30
rect 516 51 520 55
rect 539 51 542 64
rect 516 48 542 51
rect 500 22 504 26
rect 516 25 520 48
rect 717 29 721 140
rect 751 120 755 127
rect 751 119 756 120
rect 751 115 752 119
rect 759 119 763 140
rect 766 134 779 135
rect 766 130 769 134
rect 773 130 775 134
rect 766 129 779 130
rect 766 122 772 129
rect 782 123 786 140
rect 852 140 864 141
rect 868 141 948 144
rect 868 140 932 141
rect 829 129 841 135
rect 848 134 852 137
rect 936 140 948 141
rect 952 140 985 144
rect 989 140 999 144
rect 1003 140 1013 144
rect 1017 140 1023 144
rect 862 131 884 135
rect 888 131 889 135
rect 862 130 866 131
rect 848 129 852 130
rect 829 126 834 129
rect 829 125 830 126
rect 759 115 762 119
rect 766 115 767 119
rect 771 115 772 119
rect 776 115 777 119
rect 782 118 786 119
rect 821 122 830 125
rect 855 126 866 130
rect 855 122 859 126
rect 873 123 874 127
rect 878 123 889 127
rect 751 114 756 115
rect 751 106 755 114
rect 771 110 777 115
rect 758 106 759 110
rect 763 106 777 110
rect 783 108 787 111
rect 751 97 755 102
rect 751 96 756 97
rect 751 92 752 96
rect 756 92 763 95
rect 751 89 763 92
rect 767 93 771 106
rect 783 102 787 104
rect 774 98 778 102
rect 782 98 787 102
rect 774 97 787 98
rect 802 97 805 114
rect 821 108 824 122
rect 829 121 834 122
rect 838 120 859 122
rect 830 116 838 117
rect 842 118 859 120
rect 830 113 842 116
rect 830 101 834 113
rect 855 111 859 118
rect 863 116 864 120
rect 868 119 869 120
rect 868 116 880 119
rect 863 115 880 116
rect 876 112 880 115
rect 876 111 881 112
rect 844 105 850 110
rect 855 107 867 111
rect 871 107 872 111
rect 876 107 877 111
rect 844 103 846 105
rect 837 101 846 103
rect 876 106 881 107
rect 885 107 889 123
rect 876 102 880 106
rect 837 97 850 101
rect 856 98 880 102
rect 885 103 887 107
rect 830 96 834 97
rect 856 96 860 98
rect 767 89 781 93
rect 785 89 786 93
rect 843 89 844 93
rect 848 89 849 93
rect 885 94 889 103
rect 856 91 860 92
rect 865 90 866 94
rect 870 90 889 94
rect 899 92 902 131
rect 913 134 925 135
rect 913 130 918 134
rect 922 130 925 134
rect 913 129 925 130
rect 932 134 936 137
rect 946 131 968 135
rect 972 131 973 135
rect 946 130 950 131
rect 932 129 936 130
rect 913 126 918 129
rect 913 122 914 126
rect 939 126 950 130
rect 939 122 943 126
rect 957 123 958 127
rect 962 123 973 127
rect 913 121 918 122
rect 922 120 943 122
rect 914 116 922 117
rect 926 118 943 120
rect 914 113 926 116
rect 914 101 918 113
rect 939 111 943 118
rect 947 116 948 120
rect 952 119 953 120
rect 952 116 964 119
rect 947 115 964 116
rect 960 112 964 115
rect 969 116 973 123
rect 983 120 987 127
rect 983 119 988 120
rect 960 111 965 112
rect 928 105 934 110
rect 939 107 951 111
rect 955 107 956 111
rect 960 107 961 111
rect 928 103 930 105
rect 921 101 930 103
rect 960 106 965 107
rect 969 111 975 116
rect 983 115 984 119
rect 991 119 995 140
rect 998 134 1011 135
rect 998 130 1001 134
rect 1005 130 1007 134
rect 998 129 1011 130
rect 998 122 1004 129
rect 1014 123 1018 140
rect 991 115 994 119
rect 998 115 999 119
rect 1003 115 1004 119
rect 1008 115 1009 119
rect 1014 118 1018 119
rect 983 114 988 115
rect 960 102 964 106
rect 921 97 934 101
rect 940 98 964 102
rect 914 96 918 97
rect 940 96 944 98
rect 843 84 849 89
rect 927 89 928 93
rect 932 89 933 93
rect 969 94 973 111
rect 983 106 987 114
rect 1003 110 1009 115
rect 990 106 991 110
rect 995 106 1009 110
rect 940 91 944 92
rect 949 90 950 94
rect 954 90 973 94
rect 977 103 987 106
rect 977 91 980 103
rect 899 87 902 88
rect 927 84 933 89
rect 983 97 987 103
rect 983 96 988 97
rect 983 92 984 96
rect 988 92 995 95
rect 983 89 995 92
rect 999 93 1003 106
rect 1015 102 1019 105
rect 1006 98 1010 102
rect 1014 98 1019 102
rect 1006 97 1019 98
rect 999 89 1013 93
rect 1017 89 1018 93
rect 750 80 753 84
rect 757 80 763 84
rect 767 80 831 84
rect 835 80 884 84
rect 888 80 915 84
rect 919 80 968 84
rect 972 80 985 84
rect 989 80 995 84
rect 999 80 1023 84
rect 733 78 1023 80
rect 736 76 1023 78
rect 736 70 814 76
rect 840 74 884 76
rect 840 70 846 74
rect 850 70 874 74
rect 878 70 884 74
rect 844 62 850 70
rect 844 58 845 62
rect 849 58 850 62
rect 855 62 859 63
rect 864 62 870 70
rect 864 58 865 62
rect 869 58 870 62
rect 875 62 880 65
rect 879 58 880 62
rect 515 24 520 25
rect 484 18 485 22
rect 489 18 504 22
rect 507 20 515 22
rect 519 20 520 24
rect 507 18 520 20
rect 502 12 503 15
rect 480 11 503 12
rect 507 12 508 15
rect 507 11 514 12
rect 480 8 514 11
rect 518 10 524 12
rect 716 10 721 29
rect 804 30 807 56
rect 855 55 859 58
rect 875 57 880 58
rect 855 51 872 55
rect 813 29 816 42
rect 844 39 848 49
rect 852 44 857 48
rect 868 47 872 51
rect 852 36 858 40
rect 862 36 865 40
rect 852 30 856 36
rect 868 32 872 43
rect 839 27 856 30
rect 860 28 872 32
rect 876 53 880 57
rect 899 53 902 66
rect 876 50 902 53
rect 860 24 864 28
rect 876 27 880 50
rect 875 26 880 27
rect 844 20 845 24
rect 849 20 864 24
rect 867 22 875 24
rect 879 22 880 26
rect 867 20 880 22
rect 862 14 863 17
rect 518 9 721 10
rect 840 13 863 14
rect 867 14 868 17
rect 867 13 874 14
rect 840 10 874 13
rect 878 10 884 14
rect 840 9 884 10
rect 518 8 884 9
rect 480 7 884 8
rect 356 6 884 7
rect 356 5 840 6
rect 356 4 720 5
rect 356 3 480 4
rect 114 -48 117 -4
rect 673 -13 1007 -10
rect 114 -51 1009 -48
<< metal2 >>
rect 2 337 758 340
rect 762 337 853 340
rect 850 332 853 337
rect 3 324 758 327
rect 3 317 932 320
rect 3 306 705 309
rect 261 214 264 250
rect 338 189 342 286
rect 543 267 546 271
rect 390 263 533 266
rect 543 264 637 267
rect 400 244 403 263
rect 505 254 620 257
rect 399 241 403 244
rect 434 241 560 244
rect 400 215 403 241
rect 434 231 479 234
rect 476 217 479 231
rect 400 212 401 215
rect 476 214 540 217
rect 362 203 477 206
rect 362 197 365 203
rect 474 199 477 203
rect 537 199 540 214
rect 457 196 490 199
rect 338 186 404 189
rect 374 168 459 171
rect 538 171 541 195
rect 557 198 560 241
rect 561 195 594 198
rect 634 199 637 264
rect 682 265 685 297
rect 702 284 705 306
rect 702 281 838 284
rect 850 276 853 307
rect 928 290 931 317
rect 850 273 857 276
rect 903 269 906 273
rect 761 265 893 268
rect 903 266 997 269
rect 682 262 724 265
rect 650 254 710 257
rect 630 196 637 199
rect 463 168 483 171
rect 537 168 602 171
rect -16 165 307 168
rect -16 163 253 165
rect 269 163 307 165
rect 261 155 265 157
rect 261 148 264 155
rect 63 137 128 140
rect -10 129 105 132
rect 124 121 127 137
rect 206 137 291 140
rect 304 128 307 163
rect 480 154 483 168
rect 316 148 359 153
rect 480 151 542 154
rect 369 137 499 140
rect 304 124 315 128
rect -11 118 127 121
rect 28 109 35 112
rect 28 44 31 109
rect 71 110 104 113
rect 124 113 127 118
rect 175 109 208 112
rect 188 105 191 109
rect 300 105 303 111
rect 311 113 315 124
rect 369 127 373 137
rect 419 129 484 132
rect 352 123 373 127
rect 311 110 440 113
rect 480 115 483 129
rect 496 128 499 137
rect 539 133 542 151
rect 546 129 558 132
rect 496 125 534 128
rect 456 112 483 115
rect 531 116 534 125
rect 546 116 549 129
rect 562 129 647 132
rect 705 129 710 254
rect 761 217 764 265
rect 772 257 857 260
rect 817 249 918 252
rect 830 240 900 243
rect 830 217 833 240
rect 838 227 841 232
rect 838 224 901 227
rect 722 205 837 208
rect 722 199 725 205
rect 834 201 837 205
rect 898 201 901 224
rect 817 198 850 201
rect 928 200 931 256
rect 766 186 837 189
rect 734 170 819 173
rect 898 173 901 197
rect 921 197 954 200
rect 928 196 931 197
rect 994 201 997 266
rect 1005 249 1035 252
rect 1005 240 1035 243
rect 990 198 997 201
rect 823 170 843 173
rect 897 170 962 173
rect 840 156 843 170
rect 840 153 902 156
rect 729 139 859 142
rect 729 129 733 139
rect 779 131 844 134
rect 705 125 733 129
rect 531 113 549 116
rect 801 118 804 131
rect 188 102 303 105
rect 329 96 377 103
rect 264 93 265 96
rect 323 95 377 96
rect 181 70 185 93
rect 48 67 185 70
rect 262 45 265 93
rect 372 76 377 95
rect 28 41 122 44
rect 132 42 265 45
rect 345 45 349 73
rect 376 68 377 76
rect 372 67 377 68
rect 384 101 391 104
rect 280 42 349 45
rect 119 37 122 41
rect 384 36 387 101
rect 437 105 440 110
rect 427 102 460 105
rect 480 105 483 112
rect 620 111 673 114
rect 531 101 564 104
rect 544 97 547 101
rect 656 97 659 103
rect 544 94 659 97
rect 452 52 455 94
rect 539 68 542 86
rect 620 85 621 88
rect 618 37 621 85
rect 384 33 478 36
rect 488 34 631 37
rect 115 0 118 25
rect 475 29 478 33
rect 348 24 392 28
rect 453 -14 456 20
rect 670 -9 673 111
rect 689 98 737 105
rect 683 97 737 98
rect 732 78 737 97
rect 736 70 737 78
rect 732 69 737 70
rect 744 103 751 106
rect 744 38 747 103
rect 787 104 820 107
rect 840 107 843 131
rect 856 130 859 139
rect 899 135 902 153
rect 906 131 918 134
rect 856 127 894 130
rect 891 118 894 127
rect 906 118 909 131
rect 922 131 1007 134
rect 891 115 909 118
rect 979 113 1039 116
rect 813 97 816 104
rect 891 103 924 106
rect 904 99 907 103
rect 1016 99 1019 105
rect 904 96 1019 99
rect 802 62 805 93
rect 813 48 816 93
rect 899 70 902 88
rect 980 87 981 90
rect 978 39 981 87
rect 744 35 838 38
rect 848 36 991 39
rect 835 31 838 35
rect 803 24 804 25
rect 803 -3 807 24
rect -33 -19 456 -14
rect 803 -28 808 -3
rect -34 -32 808 -28
rect 814 -39 817 23
rect -32 -42 817 -39
<< ntransistor >>
rect 508 239 510 245
rect 518 239 520 245
rect 528 239 530 245
rect 735 232 737 245
rect 745 235 747 245
rect 755 238 757 252
rect 765 238 767 252
rect 785 232 787 252
rect 792 232 794 252
rect 803 232 805 246
rect 868 241 870 247
rect 878 241 880 247
rect 888 241 890 247
rect 370 208 372 217
rect 377 208 379 217
rect 389 205 391 211
rect 416 205 418 217
rect 423 205 425 217
rect 433 205 435 214
rect 443 205 445 214
rect 459 200 461 209
rect 500 205 502 217
rect 507 205 509 217
rect 517 205 519 214
rect 527 205 529 214
rect 543 200 545 209
rect 602 208 604 217
rect 609 208 611 217
rect 621 205 623 211
rect 730 210 732 219
rect 737 210 739 219
rect 749 207 751 213
rect 776 207 778 219
rect 783 207 785 219
rect 793 207 795 216
rect 803 207 805 216
rect 819 202 821 211
rect 860 207 862 219
rect 867 207 869 219
rect 877 207 879 216
rect 887 207 889 216
rect 903 202 905 211
rect 962 210 964 219
rect 969 210 971 219
rect 981 207 983 213
rect 42 97 44 103
rect 54 91 56 100
rect 61 91 63 100
rect 120 99 122 108
rect 136 94 138 103
rect 146 94 148 103
rect 156 91 158 103
rect 163 91 165 103
rect 204 99 206 108
rect 220 94 222 103
rect 230 94 232 103
rect 240 91 242 103
rect 247 91 249 103
rect 274 97 276 103
rect 286 91 288 100
rect 293 91 295 100
rect 398 89 400 95
rect 410 83 412 92
rect 417 83 419 92
rect 476 91 478 100
rect 492 86 494 95
rect 502 86 504 95
rect 39 65 41 79
rect 50 59 52 79
rect 57 59 59 79
rect 77 59 79 73
rect 87 59 89 73
rect 97 66 99 76
rect 107 66 109 79
rect 512 83 514 95
rect 519 83 521 95
rect 560 91 562 100
rect 576 86 578 95
rect 586 86 588 95
rect 596 83 598 95
rect 603 83 605 95
rect 630 89 632 95
rect 642 83 644 92
rect 649 83 651 92
rect 758 91 760 97
rect 770 85 772 94
rect 777 85 779 94
rect 836 93 838 102
rect 852 88 854 97
rect 862 88 864 97
rect 872 85 874 97
rect 879 85 881 97
rect 920 93 922 102
rect 936 88 938 97
rect 946 88 948 97
rect 956 85 958 97
rect 963 85 965 97
rect 990 91 992 97
rect 1002 85 1004 94
rect 1009 85 1011 94
rect 135 63 137 69
rect 145 63 147 69
rect 155 63 157 69
rect 491 55 493 61
rect 501 55 503 61
rect 511 55 513 61
rect 851 57 853 63
rect 861 57 863 63
rect 871 57 873 63
<< ptransistor >>
rect 508 269 510 281
rect 521 272 523 290
rect 528 272 530 290
rect 735 267 737 292
rect 748 267 750 280
rect 758 264 760 289
rect 765 264 767 289
rect 783 264 785 292
rect 793 264 795 292
rect 803 264 805 292
rect 868 271 870 283
rect 881 274 883 292
rect 888 274 890 292
rect 369 178 371 188
rect 379 178 381 188
rect 389 176 391 188
rect 415 160 417 187
rect 425 169 427 187
rect 435 169 437 187
rect 451 160 453 187
rect 499 160 501 187
rect 509 169 511 187
rect 519 169 521 187
rect 535 160 537 187
rect 601 178 603 188
rect 611 178 613 188
rect 621 176 623 188
rect 729 180 731 190
rect 739 180 741 190
rect 749 178 751 190
rect 775 162 777 189
rect 785 171 787 189
rect 795 171 797 189
rect 811 162 813 189
rect 859 162 861 189
rect 869 171 871 189
rect 879 171 881 189
rect 895 162 897 189
rect 961 180 963 190
rect 971 180 973 190
rect 981 178 983 190
rect 42 120 44 132
rect 52 120 54 130
rect 62 120 64 130
rect 128 121 130 148
rect 144 121 146 139
rect 154 121 156 139
rect 164 121 166 148
rect 212 121 214 148
rect 228 121 230 139
rect 238 121 240 139
rect 248 121 250 148
rect 274 120 276 132
rect 284 120 286 130
rect 294 120 296 130
rect 398 112 400 124
rect 408 112 410 122
rect 418 112 420 122
rect 484 113 486 140
rect 500 113 502 131
rect 510 113 512 131
rect 520 113 522 140
rect 568 113 570 140
rect 584 113 586 131
rect 594 113 596 131
rect 604 113 606 140
rect 630 112 632 124
rect 640 112 642 122
rect 650 112 652 122
rect 758 114 760 126
rect 768 114 770 124
rect 778 114 780 124
rect 844 115 846 142
rect 860 115 862 133
rect 870 115 872 133
rect 880 115 882 142
rect 928 115 930 142
rect 944 115 946 133
rect 954 115 956 133
rect 964 115 966 142
rect 990 114 992 126
rect 1000 114 1002 124
rect 1010 114 1012 124
rect 39 19 41 47
rect 49 19 51 47
rect 59 19 61 47
rect 72 19 74 47
rect 77 19 79 47
rect 84 19 86 47
rect 94 31 96 44
rect 107 19 109 44
rect 135 18 137 36
rect 142 18 144 36
rect 155 27 157 39
rect 491 10 493 28
rect 498 10 500 28
rect 511 19 513 31
rect 851 12 853 30
rect 858 12 860 30
rect 871 21 873 33
<< polycontact >>
rect 758 309 762 313
rect 519 262 523 266
rect 509 255 513 259
rect 517 254 521 258
rect 529 254 533 258
rect 742 259 746 263
rect 736 249 740 253
rect 756 256 760 260
rect 879 264 883 268
rect 775 256 779 260
rect 782 256 786 260
rect 792 256 796 260
rect 802 256 806 260
rect 869 257 873 261
rect 877 256 881 260
rect 889 256 893 260
rect 367 200 371 204
rect 447 197 451 201
rect 386 192 390 196
rect 416 191 420 195
rect 426 191 430 195
rect 531 197 535 201
rect 599 200 603 204
rect 376 168 380 172
rect 500 191 504 195
rect 510 191 514 195
rect 463 176 467 180
rect 727 202 731 206
rect 618 192 622 196
rect 807 199 811 203
rect 746 194 750 198
rect 776 193 780 197
rect 786 193 790 197
rect 891 199 895 203
rect 959 202 963 206
rect 547 176 551 180
rect 608 168 612 172
rect 736 170 740 174
rect 860 193 864 197
rect 870 193 874 197
rect 823 178 827 182
rect 978 194 982 198
rect 907 178 911 182
rect 968 170 972 174
rect 53 136 57 140
rect 114 128 118 132
rect 43 112 47 116
rect 198 128 202 132
rect 151 113 155 117
rect 161 113 165 117
rect 285 136 289 140
rect 409 128 413 132
rect 62 104 66 108
rect 130 107 134 111
rect 235 113 239 117
rect 245 113 249 117
rect 275 112 279 116
rect 214 107 218 111
rect 470 120 474 124
rect 294 104 298 108
rect 399 104 403 108
rect 554 120 558 124
rect 507 105 511 109
rect 517 105 521 109
rect 641 128 645 132
rect 769 130 773 134
rect 830 122 834 126
rect 418 96 422 100
rect 486 99 490 103
rect 591 105 595 109
rect 601 105 605 109
rect 631 104 635 108
rect 570 99 574 103
rect 759 106 763 110
rect 650 96 654 100
rect 914 122 918 126
rect 867 107 871 111
rect 877 107 881 111
rect 1001 130 1005 134
rect 778 98 782 102
rect 846 101 850 105
rect 951 107 955 111
rect 961 107 965 111
rect 991 106 995 110
rect 930 101 934 105
rect 1010 98 1014 102
rect 38 51 42 55
rect 48 51 52 55
rect 58 51 62 55
rect 65 51 69 55
rect 84 51 88 55
rect 104 58 108 62
rect 98 48 102 52
rect 132 50 136 54
rect 144 50 148 54
rect 152 49 156 53
rect 142 42 146 46
rect 488 42 492 46
rect 500 42 504 46
rect 59 -3 63 1
rect 508 41 512 45
rect 848 44 852 48
rect 860 44 864 48
rect 498 34 502 38
rect 868 43 872 47
rect 858 36 862 40
rect 83 -5 87 -1
<< ndcontact >>
rect 502 240 506 244
rect 512 240 516 244
rect 522 240 526 244
rect 532 240 536 244
rect 729 240 733 244
rect 739 236 743 240
rect 749 239 753 243
rect 759 247 763 251
rect 769 247 773 251
rect 769 240 773 244
rect 779 240 783 244
rect 796 233 800 237
rect 807 240 811 244
rect 862 242 866 246
rect 872 242 876 246
rect 882 242 886 246
rect 892 242 896 246
rect 382 218 386 222
rect 409 218 413 222
rect 364 209 368 213
rect 393 206 397 210
rect 493 218 497 222
rect 427 208 431 212
rect 437 206 441 210
rect 449 209 453 213
rect 614 218 618 222
rect 742 220 746 224
rect 769 220 773 224
rect 511 208 515 212
rect 521 206 525 210
rect 533 209 537 213
rect 596 209 600 213
rect 463 201 467 205
rect 724 211 728 215
rect 547 201 551 205
rect 625 206 629 210
rect 753 208 757 212
rect 853 220 857 224
rect 787 210 791 214
rect 797 208 801 212
rect 809 211 813 215
rect 974 220 978 224
rect 871 210 875 214
rect 881 208 885 212
rect 893 211 897 215
rect 956 211 960 215
rect 823 203 827 207
rect 907 203 911 207
rect 985 208 989 212
rect 36 98 40 102
rect 114 103 118 107
rect 198 103 202 107
rect 65 95 69 99
rect 128 95 132 99
rect 140 98 144 102
rect 150 96 154 100
rect 47 86 51 90
rect 212 95 216 99
rect 224 98 228 102
rect 234 96 238 100
rect 168 86 172 90
rect 268 98 272 102
rect 297 95 301 99
rect 252 86 256 90
rect 279 86 283 90
rect 392 90 396 94
rect 470 95 474 99
rect 554 95 558 99
rect 421 87 425 91
rect 484 87 488 91
rect 496 90 500 94
rect 506 88 510 92
rect 33 67 37 71
rect 44 74 48 78
rect 61 67 65 71
rect 71 67 75 71
rect 71 60 75 64
rect 81 60 85 64
rect 91 68 95 72
rect 101 71 105 75
rect 403 78 407 82
rect 568 87 572 91
rect 580 90 584 94
rect 590 88 594 92
rect 524 78 528 82
rect 624 90 628 94
rect 752 92 756 96
rect 830 97 834 101
rect 653 87 657 91
rect 914 97 918 101
rect 781 89 785 93
rect 844 89 848 93
rect 856 92 860 96
rect 866 90 870 94
rect 608 78 612 82
rect 635 78 639 82
rect 763 80 767 84
rect 928 89 932 93
rect 940 92 944 96
rect 950 90 954 94
rect 884 80 888 84
rect 984 92 988 96
rect 1013 89 1017 93
rect 968 80 972 84
rect 995 80 999 84
rect 111 67 115 71
rect 129 64 133 68
rect 139 64 143 68
rect 149 64 153 68
rect 159 64 163 68
rect 485 56 489 60
rect 495 56 499 60
rect 505 56 509 60
rect 515 56 519 60
rect 845 58 849 62
rect 855 58 859 62
rect 865 58 869 62
rect 875 58 879 62
<< pdcontact >>
rect 514 285 518 289
rect 502 276 506 280
rect 532 278 536 282
rect 729 275 733 279
rect 729 268 733 272
rect 740 287 744 291
rect 752 268 756 272
rect 775 287 779 291
rect 775 280 779 284
rect 787 279 791 283
rect 787 272 791 276
rect 797 287 801 291
rect 797 280 801 284
rect 874 287 878 291
rect 862 278 866 282
rect 807 272 811 276
rect 892 280 896 284
rect 807 265 811 269
rect 363 179 367 183
rect 373 183 377 187
rect 383 183 387 187
rect 393 183 397 187
rect 409 167 413 171
rect 419 175 423 179
rect 429 182 433 186
rect 445 168 449 172
rect 445 161 449 165
rect 455 182 459 186
rect 493 167 497 171
rect 503 175 507 179
rect 513 182 517 186
rect 529 168 533 172
rect 529 161 533 165
rect 539 182 543 186
rect 595 179 599 183
rect 605 183 609 187
rect 615 183 619 187
rect 625 183 629 187
rect 723 181 727 185
rect 733 185 737 189
rect 743 185 747 189
rect 753 185 757 189
rect 769 169 773 173
rect 779 177 783 181
rect 789 184 793 188
rect 805 170 809 174
rect 805 163 809 167
rect 815 184 819 188
rect 853 169 857 173
rect 863 177 867 181
rect 873 184 877 188
rect 889 170 893 174
rect 889 163 893 167
rect 899 184 903 188
rect 955 181 959 185
rect 965 185 969 189
rect 975 185 979 189
rect 985 185 989 189
rect 36 121 40 125
rect 46 121 50 125
rect 56 121 60 125
rect 66 125 70 129
rect 122 122 126 126
rect 132 143 136 147
rect 132 136 136 140
rect 148 122 152 126
rect 158 129 162 133
rect 168 137 172 141
rect 206 122 210 126
rect 216 143 220 147
rect 216 136 220 140
rect 232 122 236 126
rect 242 129 246 133
rect 252 137 256 141
rect 268 121 272 125
rect 278 121 282 125
rect 288 121 292 125
rect 298 125 302 129
rect 392 113 396 117
rect 402 113 406 117
rect 412 113 416 117
rect 422 117 426 121
rect 478 114 482 118
rect 488 135 492 139
rect 488 128 492 132
rect 504 114 508 118
rect 514 121 518 125
rect 524 129 528 133
rect 562 114 566 118
rect 572 135 576 139
rect 572 128 576 132
rect 588 114 592 118
rect 598 121 602 125
rect 608 129 612 133
rect 624 113 628 117
rect 634 113 638 117
rect 644 113 648 117
rect 654 117 658 121
rect 752 115 756 119
rect 762 115 766 119
rect 772 115 776 119
rect 782 119 786 123
rect 838 116 842 120
rect 848 137 852 141
rect 848 130 852 134
rect 864 116 868 120
rect 874 123 878 127
rect 884 131 888 135
rect 922 116 926 120
rect 932 137 936 141
rect 932 130 936 134
rect 948 116 952 120
rect 958 123 962 127
rect 968 131 972 135
rect 984 115 988 119
rect 994 115 998 119
rect 1004 115 1008 119
rect 1014 119 1018 123
rect 33 42 37 46
rect 33 35 37 39
rect 43 27 47 31
rect 43 20 47 24
rect 53 35 57 39
rect 53 28 57 32
rect 65 27 69 31
rect 65 20 69 24
rect 88 39 92 43
rect 100 20 104 24
rect 111 39 115 43
rect 111 32 115 36
rect 129 26 133 30
rect 159 28 163 32
rect 147 19 151 23
rect 485 18 489 22
rect 515 20 519 24
rect 845 20 849 24
rect 503 11 507 15
rect 875 22 879 26
rect 863 13 867 17
<< m2contact >>
rect 681 344 685 348
rect 758 336 762 340
rect 849 328 853 332
rect 758 324 762 328
rect 850 307 854 311
rect 681 297 685 301
rect 338 286 342 290
rect 260 250 264 254
rect 501 254 505 258
rect 542 271 546 275
rect 927 286 931 290
rect 838 280 842 284
rect 533 263 537 267
rect 620 254 624 258
rect 646 254 650 258
rect 429 241 434 245
rect 430 231 434 235
rect 260 210 264 214
rect 261 157 265 161
rect 59 136 63 140
rect 105 128 109 132
rect 35 108 39 112
rect 67 110 71 114
rect 104 110 108 114
rect 124 109 128 113
rect 171 109 175 113
rect 202 136 206 140
rect 260 144 264 148
rect 311 148 316 153
rect 291 136 295 140
rect 208 109 212 113
rect 181 93 185 97
rect 260 93 264 97
rect 299 111 303 115
rect 362 193 366 197
rect 401 211 405 215
rect 370 168 374 172
rect 404 186 408 190
rect 453 195 457 199
rect 490 195 494 199
rect 537 195 541 199
rect 557 194 561 198
rect 594 194 598 198
rect 626 196 630 200
rect 459 168 463 172
rect 602 168 606 172
rect 724 261 728 265
rect 768 256 772 260
rect 813 249 817 253
rect 857 272 861 276
rect 857 257 861 261
rect 902 273 906 277
rect 893 265 897 269
rect 927 256 931 260
rect 918 249 922 253
rect 1001 249 1005 253
rect 837 232 841 236
rect 900 240 904 244
rect 1001 240 1005 244
rect 359 148 365 154
rect 323 96 329 103
rect 345 123 352 129
rect 44 67 48 71
rect 128 41 132 45
rect 119 33 123 37
rect 275 42 280 46
rect 115 25 119 29
rect 342 73 350 80
rect 343 24 348 30
rect 415 128 419 132
rect 538 129 542 133
rect 451 112 456 118
rect 391 100 395 104
rect 423 102 427 106
rect 460 102 464 106
rect 451 94 455 98
rect 480 101 484 105
rect 527 101 531 105
rect 558 128 562 132
rect 616 111 620 115
rect 647 128 651 132
rect 564 101 568 105
rect 539 86 543 90
rect 616 85 620 89
rect 655 103 659 107
rect 722 195 726 199
rect 761 213 765 217
rect 830 213 836 217
rect 813 197 817 201
rect 730 170 734 174
rect 762 185 766 189
rect 850 197 854 201
rect 837 186 841 190
rect 897 197 901 201
rect 917 196 921 200
rect 954 196 958 200
rect 986 198 990 202
rect 819 170 823 174
rect 962 170 966 174
rect 683 98 689 105
rect 368 68 376 76
rect 538 64 542 68
rect 451 47 456 52
rect 392 22 398 28
rect 484 33 488 37
rect 452 20 457 26
rect 475 25 479 29
rect 775 130 779 134
rect 898 131 902 135
rect 801 114 805 118
rect 751 102 755 106
rect 783 104 787 108
rect 820 104 824 108
rect 840 103 844 107
rect 887 103 891 107
rect 802 93 806 97
rect 812 93 816 97
rect 918 130 922 134
rect 924 103 928 107
rect 975 111 979 116
rect 1007 130 1011 134
rect 899 88 903 92
rect 976 87 980 91
rect 1015 105 1019 109
rect 728 70 736 78
rect 802 56 807 62
rect 898 66 902 70
rect 812 42 817 48
rect 804 24 809 30
rect 844 35 848 39
rect 813 23 818 29
rect 835 27 839 31
rect 114 -4 118 0
rect 669 -13 673 -9
<< psubstratepcontact >>
rect 503 228 507 232
rect 531 228 535 232
rect 863 230 867 234
rect 891 230 895 234
rect 392 218 396 222
rect 462 218 466 222
rect 546 218 550 222
rect 624 218 628 222
rect 752 220 756 224
rect 822 220 826 224
rect 906 220 910 224
rect 984 220 988 224
rect 37 86 41 90
rect 115 86 119 90
rect 199 86 203 90
rect 269 86 273 90
rect 130 76 134 80
rect 158 76 162 80
rect 393 78 397 82
rect 471 78 475 82
rect 555 78 559 82
rect 625 78 629 82
rect 753 80 757 84
rect 831 80 835 84
rect 915 80 919 84
rect 985 80 989 84
rect 486 68 490 72
rect 514 68 518 72
rect 846 70 850 74
rect 874 70 878 74
<< nsubstratencontact >>
rect 503 288 507 292
rect 863 290 867 294
rect 364 158 368 162
rect 378 158 382 162
rect 392 158 396 162
rect 429 158 433 162
rect 513 158 517 162
rect 596 158 600 162
rect 610 158 614 162
rect 624 158 628 162
rect 724 160 728 164
rect 738 160 742 164
rect 752 160 756 164
rect 789 160 793 164
rect 873 160 877 164
rect 956 160 960 164
rect 970 160 974 164
rect 984 160 988 164
rect 37 146 41 150
rect 51 146 55 150
rect 65 146 69 150
rect 148 146 152 150
rect 232 146 236 150
rect 269 146 273 150
rect 283 146 287 150
rect 297 146 301 150
rect 393 138 397 142
rect 407 138 411 142
rect 421 138 425 142
rect 504 138 508 142
rect 588 138 592 142
rect 625 138 629 142
rect 639 138 643 142
rect 653 138 657 142
rect 753 140 757 144
rect 767 140 771 144
rect 781 140 785 144
rect 864 140 868 144
rect 948 140 952 144
rect 985 140 989 144
rect 999 140 1003 144
rect 1013 140 1017 144
rect 158 16 162 20
rect 514 8 518 12
rect 874 10 878 14
<< psubstratepdiff >>
rect 502 232 536 233
rect 502 228 503 232
rect 507 228 531 232
rect 535 228 536 232
rect 862 234 896 235
rect 862 230 863 234
rect 867 230 891 234
rect 895 230 896 234
rect 862 229 896 230
rect 502 227 536 228
rect 391 222 397 223
rect 391 218 392 222
rect 396 218 397 222
rect 391 217 397 218
rect 461 222 467 223
rect 461 218 462 222
rect 466 218 467 222
rect 461 217 467 218
rect 545 222 551 223
rect 545 218 546 222
rect 550 218 551 222
rect 545 217 551 218
rect 623 222 629 223
rect 623 218 624 222
rect 628 218 629 222
rect 751 224 757 225
rect 751 220 752 224
rect 756 220 757 224
rect 751 219 757 220
rect 623 217 629 218
rect 821 224 827 225
rect 821 220 822 224
rect 826 220 827 224
rect 821 219 827 220
rect 905 224 911 225
rect 905 220 906 224
rect 910 220 911 224
rect 905 219 911 220
rect 983 224 989 225
rect 983 220 984 224
rect 988 220 989 224
rect 983 219 989 220
rect 36 90 42 91
rect 36 86 37 90
rect 41 86 42 90
rect 36 85 42 86
rect 114 90 120 91
rect 114 86 115 90
rect 119 86 120 90
rect 114 85 120 86
rect 198 90 204 91
rect 198 86 199 90
rect 203 86 204 90
rect 198 85 204 86
rect 268 90 274 91
rect 268 86 269 90
rect 273 86 274 90
rect 268 85 274 86
rect 392 82 398 83
rect 129 80 163 81
rect 129 76 130 80
rect 134 76 158 80
rect 162 76 163 80
rect 392 78 393 82
rect 397 78 398 82
rect 392 77 398 78
rect 470 82 476 83
rect 470 78 471 82
rect 475 78 476 82
rect 470 77 476 78
rect 554 82 560 83
rect 554 78 555 82
rect 559 78 560 82
rect 554 77 560 78
rect 752 84 758 85
rect 624 82 630 83
rect 624 78 625 82
rect 629 78 630 82
rect 624 77 630 78
rect 752 80 753 84
rect 757 80 758 84
rect 752 79 758 80
rect 830 84 836 85
rect 830 80 831 84
rect 835 80 836 84
rect 830 79 836 80
rect 914 84 920 85
rect 914 80 915 84
rect 919 80 920 84
rect 914 79 920 80
rect 984 84 990 85
rect 984 80 985 84
rect 989 80 990 84
rect 984 79 990 80
rect 129 75 163 76
rect 845 74 879 75
rect 485 72 519 73
rect 485 68 486 72
rect 490 68 514 72
rect 518 68 519 72
rect 845 70 846 74
rect 850 70 874 74
rect 878 70 879 74
rect 845 69 879 70
rect 485 67 519 68
<< nsubstratendiff >>
rect 502 292 508 293
rect 502 288 503 292
rect 507 288 508 292
rect 502 287 508 288
rect 862 294 868 295
rect 862 290 863 294
rect 867 290 868 294
rect 862 289 868 290
rect 363 162 397 163
rect 363 158 364 162
rect 368 158 378 162
rect 382 158 392 162
rect 396 158 397 162
rect 428 162 434 163
rect 363 157 397 158
rect 428 158 429 162
rect 433 158 434 162
rect 512 162 518 163
rect 428 157 434 158
rect 512 158 513 162
rect 517 158 518 162
rect 723 164 757 165
rect 595 162 629 163
rect 512 157 518 158
rect 595 158 596 162
rect 600 158 610 162
rect 614 158 624 162
rect 628 158 629 162
rect 723 160 724 164
rect 728 160 738 164
rect 742 160 752 164
rect 756 160 757 164
rect 788 164 794 165
rect 723 159 757 160
rect 788 160 789 164
rect 793 160 794 164
rect 872 164 878 165
rect 788 159 794 160
rect 872 160 873 164
rect 877 160 878 164
rect 955 164 989 165
rect 872 159 878 160
rect 955 160 956 164
rect 960 160 970 164
rect 974 160 984 164
rect 988 160 989 164
rect 955 159 989 160
rect 595 157 629 158
rect 36 150 70 151
rect 36 146 37 150
rect 41 146 51 150
rect 55 146 65 150
rect 69 146 70 150
rect 147 150 153 151
rect 36 145 70 146
rect 147 146 148 150
rect 152 146 153 150
rect 231 150 237 151
rect 147 145 153 146
rect 231 146 232 150
rect 236 146 237 150
rect 268 150 302 151
rect 231 145 237 146
rect 268 146 269 150
rect 273 146 283 150
rect 287 146 297 150
rect 301 146 302 150
rect 268 145 302 146
rect 752 144 786 145
rect 392 142 426 143
rect 392 138 393 142
rect 397 138 407 142
rect 411 138 421 142
rect 425 138 426 142
rect 503 142 509 143
rect 392 137 426 138
rect 503 138 504 142
rect 508 138 509 142
rect 587 142 593 143
rect 503 137 509 138
rect 587 138 588 142
rect 592 138 593 142
rect 624 142 658 143
rect 587 137 593 138
rect 624 138 625 142
rect 629 138 639 142
rect 643 138 653 142
rect 657 138 658 142
rect 752 140 753 144
rect 757 140 767 144
rect 771 140 781 144
rect 785 140 786 144
rect 863 144 869 145
rect 752 139 786 140
rect 624 137 658 138
rect 863 140 864 144
rect 868 140 869 144
rect 947 144 953 145
rect 863 139 869 140
rect 947 140 948 144
rect 952 140 953 144
rect 984 144 1018 145
rect 947 139 953 140
rect 984 140 985 144
rect 989 140 999 144
rect 1003 140 1013 144
rect 1017 140 1018 144
rect 984 139 1018 140
rect 157 20 163 21
rect 157 16 158 20
rect 162 16 163 20
rect 157 15 163 16
rect 513 12 519 13
rect 873 14 879 15
rect 513 8 514 12
rect 518 8 519 12
rect 873 10 874 14
rect 878 10 879 14
rect 873 9 879 10
rect 513 7 519 8
<< labels >>
rlabel metal1 143 86 143 86 6 vss
rlabel metal1 143 150 143 150 6 vdd
rlabel metal1 227 86 227 86 6 vss
rlabel metal1 227 150 227 150 6 vdd
rlabel metal1 53 86 53 86 6 vss
rlabel metal1 53 150 53 150 6 vdd
rlabel metal1 285 150 285 150 6 vdd
rlabel metal1 285 86 285 86 6 vss
rlabel metal1 146 80 146 80 2 vss
rlabel metal1 146 16 146 16 2 vdd
rlabel metal1 70 17 70 17 2 vdd
rlabel metal1 70 81 70 81 2 vss
rlabel metal1 502 8 502 8 2 vdd
rlabel metal1 641 142 641 142 6 vdd
rlabel metal1 409 142 409 142 6 vdd
rlabel metal1 583 142 583 142 6 vdd
rlabel metal1 499 142 499 142 6 vdd
rlabel metal1 499 78 499 78 6 vss
rlabel metal1 519 292 519 292 6 vdd
rlabel metal1 519 228 519 228 6 vss
rlabel metal1 380 222 380 222 2 vss
rlabel metal1 380 158 380 158 2 vdd
rlabel metal1 612 158 612 158 2 vdd
rlabel metal1 612 222 612 222 2 vss
rlabel metal1 438 158 438 158 2 vdd
rlabel metal1 522 158 522 158 2 vdd
rlabel metal1 862 10 862 10 2 vdd
rlabel metal1 1001 144 1001 144 6 vdd
rlabel metal1 769 144 769 144 6 vdd
rlabel metal1 943 144 943 144 6 vdd
rlabel metal1 859 144 859 144 6 vdd
rlabel metal1 859 80 859 80 6 vss
rlabel metal1 879 294 879 294 6 vdd
rlabel metal1 879 230 879 230 6 vss
rlabel metal1 740 224 740 224 2 vss
rlabel metal1 740 160 740 160 2 vdd
rlabel metal1 972 160 972 160 2 vdd
rlabel metal1 972 224 972 224 2 vss
rlabel metal1 798 160 798 160 2 vdd
rlabel metal1 882 160 882 160 2 vdd
rlabel metal1 511 260 511 260 1 cout3_n_A2
rlabel m2contact 503 256 503 256 1 c3_A2
rlabel metal1 863 258 863 258 1 c5_A2
rlabel metal1 871 262 871 262 1 cout5_n_A2
rlabel metal1 980 212 980 212 1 n18_A2
rlabel metal1 967 192 967 192 1 n18_n_A2
rlabel polycontact 894 200 894 200 1 a5_A2
rlabel metal1 910 176 910 176 1 b5_A2
rlabel metal1 878 195 878 195 1 b5_n_A2
rlabel polycontact 863 195 863 195 1 a5_n_A2
rlabel metal1 854 192 854 192 1 xor_5_A2
rlabel m2contact 820 172 820 172 1 c4_A2
rlabel metal1 798 176 798 176 1 n20_A2
rlabel metal1 770 192 770 192 1 s6_A2
rlabel polycontact 778 194 778 194 1 n19_A2
rlabel metal1 756 196 756 196 1 n21_A2
rlabel metal1 742 196 742 196 1 zc5_n_A2
rlabel metal1 620 210 620 210 1 n10_A2
rlabel metal1 607 190 607 190 1 n1_n_A2
rlabel metal1 518 193 518 193 1 b3n_A2
rlabel polycontact 503 193 503 193 1 a3n_A2
rlabel metal1 494 190 494 190 1 xor_3_A2
rlabel metal2 458 170 458 170 1 c2_A2
rlabel metal1 438 174 438 174 1 n12_A2
rlabel metal1 410 190 410 190 1 s4_A2
rlabel ntransistor 417 207 417 207 1 n11_A2
rlabel metal1 396 194 396 194 1 n13_A2
rlabel metal1 382 194 382 194 1 zc3_n_A2
rlabel metal1 999 108 999 108 1 zc4_n_A2
rlabel metal1 985 108 985 108 1 n16_A2
rlabel metal1 971 112 971 112 1 s5_A2
rlabel metal1 948 129 948 129 1 n14_A2
rlabel metal2 907 132 907 132 1 c3_A2
rlabel metal1 887 112 887 112 1 xor_4_A2
rlabel ptransistor 871 117 871 117 1 a4n_A2
rlabel metal1 839 100 839 100 1 a4_A2
rlabel metal1 832 106 832 106 1 b4n_A2
rlabel metal1 831 129 831 129 1 b4_A2
rlabel metal1 774 112 774 112 1 n17_n_A2
rlabel metal1 761 92 761 92 1 n17_A2
rlabel metal2 712 127 712 127 1 c3_A2
rlabel metal1 639 106 639 106 1 zc2_n_A2
rlabel metal1 625 106 625 106 1 n8_A2
rlabel metal1 611 110 611 110 1 s3_A2
rlabel metal1 588 127 588 127 1 n6_A2
rlabel metal2 547 130 547 130 1 s2_A2
rlabel metal1 527 110 527 110 1 xor_2_A2
rlabel ptransistor 511 115 511 115 1 a2n_A2
rlabel metal1 479 98 479 98 1 a2_A2
rlabel metal1 472 104 472 104 1 b2n_A2
rlabel metal1 471 127 471 127 1 b2_A2
rlabel metal1 401 90 401 90 1 n9_A2
rlabel m2contact 349 126 349 126 1 s2_A2
rlabel metal1 283 114 283 114 1 zc1_n_A2
rlabel metal1 269 114 269 114 1 c1_A2
rlabel metal1 255 118 255 118 1 s1_A2
rlabel metal1 231 133 231 133 1 n3_A2
rlabel metal1 171 118 171 118 1 xor1_A2
rlabel metal1 159 139 159 139 1 bn_A2
rlabel ndcontact 141 100 141 100 1 a1n_A2
rlabel polycontact 131 110 131 110 1 a1_A2
rlabel metal1 116 112 116 112 1 b1n_A2
rlabel polycontact 115 130 115 130 1 b1_A2
rlabel metal1 45 98 45 98 1 n5_A2
rlabel ndcontact 34 69 34 69 1 co_A2
rlabel polycontact 40 53 40 53 1 con_A2
rlabel polycontact 60 53 60 53 1 a_A2
rlabel metal1 73 66 73 66 1 n2_A2
rlabel ntransistor 88 62 88 62 1 son_A2
rlabel polycontact 100 50 100 50 1 con_A2
rlabel metal1 82 49 82 49 1 b_A2
rlabel metal1 114 53 114 53 1 so_A2
rlabel metal1 162 52 162 52 1 s2_A2
rlabel metal1 518 44 518 44 1 c2_A2
rlabel metal1 510 40 510 40 1 cout2_n_A2
rlabel metal1 870 42 870 42 1 cout4_n_A2
rlabel metal1 878 46 878 46 1 c4_A2
rlabel metal1 154 48 154 48 1 cout_n_A2
rlabel polycontact 533 199 533 199 1 a3_A2
rlabel metal1 550 174 550 174 1 b3_A2
rlabel polycontact 963 109 963 109 1 n15_A2
rlabel polycontact 603 107 603 107 1 n7_A2
rlabel polycontact 247 115 247 115 1 n4_A2
rlabel metal1 774 230 774 230 6 vss
rlabel metal1 774 294 774 294 6 vdd
rlabel polycontact 758 257 758 257 1 c5_A1
rlabel metal1 810 253 810 253 1 s8_A2
rlabel metal1 771 245 771 245 1 n2_7_A2
rlabel ptransistor 784 274 784 274 1 s8_n_A2
rlabel polycontact 738 251 738 251 1 s7_n_A2
rlabel metal1 730 258 730 258 1 s7_A2
rlabel metal1 58 116 58 116 1 n1_A2
rlabel metal2 -8 120 -8 120 1 a1_A2
rlabel metal2 -6 130 -6 130 1 b1_A2
rlabel metal1 414 107 414 107 1 n9_n_A2
rlabel metal2 -8 166 -8 166 1 b2_A2
rlabel metal2 -28 -19 -28 -19 2 a2_A2
rlabel metal2 -28 -41 -28 -41 1 b4_A2
rlabel metal2 -26 -31 -26 -31 1 a4_A2
rlabel metal1 8 233 8 233 1 a3_A2
rlabel metal1 7 242 7 242 1 b3_A2
rlabel metal2 6 308 6 308 5 a5_A2
rlabel metal2 5 319 5 319 5 b5_A2
rlabel metal2 1032 251 1032 251 7 s8_A2
rlabel metal1 1054 346 1054 346 5 s7_A2
rlabel metal1 1056 362 1056 362 6 s4_A2
rlabel metal1 1051 379 1051 379 5 s1_A2
rlabel metal1 1005 -12 1005 -12 1 s3_A2
rlabel metal2 1033 115 1033 115 1 s5_A2
rlabel metal1 1007 -49 1007 -49 1 so_A2
rlabel metal2 1032 242 1032 242 1 s6_A2
rlabel metal2 4 339 4 339 1 c5_A2
rlabel metal2 5 326 5 326 1 c5_A1
rlabel polycontact 85 -3 85 -3 2 b_A2
rlabel polycontact 61 -1 61 -1 3 a_A2
<< end >>
