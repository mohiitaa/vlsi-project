magic
tech scmos
timestamp 1520243457
<< nwell >>
rect -17 4 -5 15
rect 5 4 17 15
<< polysilicon >>
rect -12 11 -10 13
rect 10 11 12 13
rect -12 3 -10 8
rect -11 -1 -10 3
rect -12 -5 -10 -1
rect 10 3 12 8
rect 10 -1 11 3
rect 10 -5 12 -1
rect -12 -10 -10 -8
rect 10 -10 12 -8
<< ndiffusion >>
rect -13 -8 -12 -5
rect -10 -8 -9 -5
rect 9 -8 10 -5
rect 12 -8 13 -5
<< pdiffusion >>
rect -13 8 -12 11
rect -10 8 -9 11
rect 9 8 10 11
rect 12 8 13 11
<< metal1 >>
rect -17 17 17 20
rect -17 12 -14 17
rect 14 12 17 17
rect -8 3 -5 8
rect -2 8 5 11
rect -2 3 1 8
rect -8 0 1 3
rect -8 -4 -5 0
rect -17 -11 -14 -8
rect 5 -11 8 -8
rect -17 -14 8 -11
rect 14 -19 17 -8
rect -17 -22 17 -19
<< ntransistor >>
rect -12 -8 -10 -5
rect 10 -8 12 -5
<< ptransistor >>
rect -12 8 -10 11
rect 10 8 12 11
<< polycontact >>
rect -15 -1 -11 3
rect 11 -1 15 3
<< ndcontact >>
rect -17 -8 -13 -4
rect -9 -8 -5 -4
rect 5 -8 9 -4
rect 13 -8 17 -4
<< pdcontact >>
rect -17 8 -13 12
rect -9 8 -5 12
rect 5 8 9 12
rect 13 8 17 12
<< labels >>
rlabel polycontact -13 1 -13 1 3 A
rlabel polycontact 13 1 13 1 7 B
rlabel metal1 -1 19 -1 19 5 vdd
rlabel metal1 0 -21 0 -21 1 gnd
rlabel metal1 0 2 0 2 1 out
<< end >>
