magic
tech scmos
timestamp 1523031569
<< nwell >>
rect 3 116 182 142
rect 195 116 236 142
rect 251 116 292 142
rect 305 116 346 142
rect 99 11 186 37
rect 199 11 240 37
rect 255 11 296 37
rect 309 11 350 37
<< polysilicon >>
rect 40 129 42 131
rect 112 129 114 135
rect 151 129 153 135
rect 172 129 174 135
rect 205 129 207 135
rect 226 129 228 135
rect 261 129 263 135
rect 282 129 284 135
rect 315 129 317 135
rect 336 129 338 135
rect 40 112 42 123
rect 112 111 114 123
rect 151 111 153 123
rect 172 111 174 123
rect 205 111 207 123
rect 226 111 228 123
rect 261 111 263 123
rect 282 111 284 123
rect 315 111 317 123
rect 336 111 338 123
rect 40 90 42 108
rect 152 107 153 111
rect 173 107 174 111
rect 206 107 207 111
rect 227 107 228 111
rect 262 107 263 111
rect 283 107 284 111
rect 316 107 317 111
rect 337 107 338 111
rect 40 84 42 87
rect 112 89 114 107
rect 151 92 153 107
rect 172 92 174 107
rect 205 92 207 107
rect 226 92 228 107
rect 261 92 263 107
rect 282 92 284 107
rect 315 92 317 107
rect 336 92 338 107
rect 112 83 114 86
rect 151 83 153 86
rect 172 83 174 86
rect 205 83 207 86
rect 226 83 228 86
rect 261 83 263 86
rect 282 83 284 86
rect 315 83 317 86
rect 336 83 338 86
rect 116 67 118 70
rect 155 67 157 70
rect 176 67 178 70
rect 209 67 211 70
rect 230 67 232 70
rect 265 67 267 70
rect 286 67 288 70
rect 319 67 321 70
rect 340 67 342 70
rect 116 46 118 64
rect 155 46 157 61
rect 176 46 178 61
rect 209 46 211 61
rect 230 46 232 61
rect 265 46 267 61
rect 286 46 288 61
rect 319 46 321 61
rect 340 46 342 61
rect 156 42 157 46
rect 177 42 178 46
rect 210 42 211 46
rect 231 42 232 46
rect 266 42 267 46
rect 287 42 288 46
rect 320 42 321 46
rect 341 42 342 46
rect 116 30 118 42
rect 155 30 157 42
rect 176 30 178 42
rect 209 30 211 42
rect 230 30 232 42
rect 265 30 267 42
rect 286 30 288 42
rect 319 30 321 42
rect 340 30 342 42
rect 116 18 118 24
rect 155 18 157 24
rect 176 18 178 24
rect 209 18 211 24
rect 230 18 232 24
rect 265 18 267 24
rect 286 18 288 24
rect 319 18 321 24
rect 340 18 342 24
<< ndiffusion >>
rect 29 87 40 90
rect 42 87 59 90
rect 141 91 151 92
rect 101 86 112 89
rect 114 86 131 89
rect 141 87 143 91
rect 147 87 151 91
rect 141 86 151 87
rect 153 86 172 92
rect 174 91 182 92
rect 174 87 177 91
rect 181 87 182 91
rect 174 86 182 87
rect 195 91 205 92
rect 195 87 197 91
rect 201 87 205 91
rect 195 86 205 87
rect 207 86 226 92
rect 228 91 236 92
rect 228 87 231 91
rect 235 87 236 91
rect 228 86 236 87
rect 251 91 261 92
rect 251 87 253 91
rect 257 87 261 91
rect 251 86 261 87
rect 263 86 282 92
rect 284 91 292 92
rect 284 87 287 91
rect 291 87 292 91
rect 284 86 292 87
rect 305 91 315 92
rect 305 87 307 91
rect 311 87 315 91
rect 305 86 315 87
rect 317 86 336 92
rect 338 91 346 92
rect 338 87 341 91
rect 345 87 346 91
rect 338 86 346 87
rect 105 64 116 67
rect 118 64 135 67
rect 145 66 155 67
rect 145 62 147 66
rect 151 62 155 66
rect 145 61 155 62
rect 157 61 176 67
rect 178 66 186 67
rect 178 62 181 66
rect 185 62 186 66
rect 178 61 186 62
rect 199 66 209 67
rect 199 62 201 66
rect 205 62 209 66
rect 199 61 209 62
rect 211 61 230 67
rect 232 66 240 67
rect 232 62 235 66
rect 239 62 240 66
rect 232 61 240 62
rect 255 66 265 67
rect 255 62 257 66
rect 261 62 265 66
rect 255 61 265 62
rect 267 61 286 67
rect 288 66 296 67
rect 288 62 291 66
rect 295 62 296 66
rect 288 61 296 62
rect 309 66 319 67
rect 309 62 311 66
rect 315 62 319 66
rect 309 61 319 62
rect 321 61 340 67
rect 342 66 350 67
rect 342 62 345 66
rect 349 62 350 66
rect 342 61 350 62
<< pdiffusion >>
rect 9 128 40 129
rect 9 124 14 128
rect 18 124 40 128
rect 9 123 40 124
rect 42 124 58 129
rect 64 124 77 129
rect 42 123 77 124
rect 97 128 112 129
rect 101 124 112 128
rect 97 123 112 124
rect 114 128 134 129
rect 114 124 130 128
rect 114 123 134 124
rect 141 128 151 129
rect 141 124 143 128
rect 147 124 151 128
rect 141 123 151 124
rect 153 128 172 129
rect 153 124 160 128
rect 164 124 172 128
rect 153 123 172 124
rect 174 128 182 129
rect 174 124 177 128
rect 181 124 182 128
rect 174 123 182 124
rect 195 128 205 129
rect 195 124 197 128
rect 201 124 205 128
rect 195 123 205 124
rect 207 128 226 129
rect 207 124 214 128
rect 218 124 226 128
rect 207 123 226 124
rect 228 128 236 129
rect 228 124 231 128
rect 235 124 236 128
rect 228 123 236 124
rect 251 128 261 129
rect 251 124 253 128
rect 257 124 261 128
rect 251 123 261 124
rect 263 128 282 129
rect 263 124 270 128
rect 274 124 282 128
rect 263 123 282 124
rect 284 128 292 129
rect 284 124 287 128
rect 291 124 292 128
rect 284 123 292 124
rect 305 128 315 129
rect 305 124 307 128
rect 311 124 315 128
rect 305 123 315 124
rect 317 128 336 129
rect 317 124 324 128
rect 328 124 336 128
rect 317 123 336 124
rect 338 128 346 129
rect 338 124 341 128
rect 345 124 346 128
rect 338 123 346 124
rect 101 29 116 30
rect 105 25 116 29
rect 101 24 116 25
rect 118 29 138 30
rect 118 25 134 29
rect 118 24 138 25
rect 145 29 155 30
rect 145 25 147 29
rect 151 25 155 29
rect 145 24 155 25
rect 157 29 176 30
rect 157 25 164 29
rect 168 25 176 29
rect 157 24 176 25
rect 178 29 186 30
rect 178 25 181 29
rect 185 25 186 29
rect 178 24 186 25
rect 199 29 209 30
rect 199 25 201 29
rect 205 25 209 29
rect 199 24 209 25
rect 211 29 230 30
rect 211 25 218 29
rect 222 25 230 29
rect 211 24 230 25
rect 232 29 240 30
rect 232 25 235 29
rect 239 25 240 29
rect 232 24 240 25
rect 255 29 265 30
rect 255 25 257 29
rect 261 25 265 29
rect 255 24 265 25
rect 267 29 286 30
rect 267 25 274 29
rect 278 25 286 29
rect 267 24 286 25
rect 288 29 296 30
rect 288 25 291 29
rect 295 25 296 29
rect 288 24 296 25
rect 309 29 319 30
rect 309 25 311 29
rect 315 25 319 29
rect 309 24 319 25
rect 321 29 340 30
rect 321 25 328 29
rect 332 25 340 29
rect 321 24 340 25
rect 342 29 350 30
rect 342 25 345 29
rect 349 25 350 29
rect 342 24 350 25
<< metal1 >>
rect -2 147 364 150
rect 14 128 17 147
rect 59 130 63 132
rect 97 128 100 147
rect 160 128 163 147
rect 170 142 173 147
rect 214 128 217 147
rect 224 142 227 147
rect 270 128 273 147
rect 280 142 283 147
rect 324 128 327 147
rect 334 142 337 147
rect 59 113 63 124
rect 42 109 45 112
rect 59 103 62 113
rect 114 108 117 111
rect 59 99 60 103
rect 131 102 134 124
rect 144 119 147 124
rect 177 119 180 124
rect 144 116 180 119
rect 146 108 148 111
rect 168 108 169 111
rect 177 107 180 116
rect 198 119 201 124
rect 231 119 234 124
rect 198 116 234 119
rect 254 119 257 124
rect 287 119 290 124
rect 254 116 290 119
rect 308 119 311 124
rect 341 119 344 124
rect 308 116 344 119
rect 184 107 187 116
rect 198 111 205 112
rect 198 109 202 111
rect 219 107 223 110
rect 177 104 187 107
rect 59 91 62 99
rect 131 98 132 102
rect 131 90 134 98
rect 177 91 180 104
rect 219 103 222 107
rect 231 104 234 116
rect 287 115 290 116
rect 255 108 258 111
rect 231 101 250 104
rect 231 91 234 101
rect 279 105 282 107
rect 267 97 270 103
rect 281 101 282 105
rect 279 100 282 101
rect 244 94 270 97
rect 287 91 290 111
rect 311 107 312 110
rect 330 111 336 112
rect 330 109 333 111
rect 311 98 314 107
rect 341 106 344 116
rect 313 94 314 98
rect 341 91 344 102
rect 25 81 28 87
rect 97 81 100 86
rect 143 81 146 87
rect 197 81 200 87
rect 253 81 256 87
rect 307 81 310 87
rect 1 78 346 81
rect 169 75 174 78
rect 275 75 279 78
rect 101 72 350 75
rect 101 67 104 72
rect 147 66 150 72
rect 201 66 204 72
rect 257 66 260 72
rect 311 66 314 72
rect 135 55 138 63
rect 135 51 136 55
rect 118 42 121 45
rect 135 29 138 51
rect 181 49 184 62
rect 181 46 191 49
rect 223 46 226 50
rect 235 52 238 62
rect 235 49 254 52
rect 283 52 286 53
rect 150 42 152 45
rect 172 42 173 45
rect 181 37 184 46
rect 148 34 184 37
rect 148 29 151 34
rect 181 29 184 34
rect 188 37 191 46
rect 202 42 206 44
rect 223 43 227 46
rect 202 41 209 42
rect 235 37 238 49
rect 285 48 286 52
rect 283 46 286 48
rect 259 42 262 45
rect 291 42 294 62
rect 317 55 318 59
rect 315 46 318 55
rect 345 51 348 62
rect 315 43 316 46
rect 334 42 337 44
rect 334 41 340 42
rect 291 37 294 38
rect 345 37 348 47
rect 202 34 238 37
rect 202 29 205 34
rect 235 29 238 34
rect 258 34 294 37
rect 258 29 261 34
rect 291 29 294 34
rect 312 34 348 37
rect 312 29 315 34
rect 345 29 348 34
rect 101 6 104 25
rect 164 6 167 25
rect 174 6 177 11
rect 218 6 221 25
rect 228 6 231 11
rect 274 6 277 25
rect 284 6 287 11
rect 328 6 331 25
rect 338 6 341 11
rect 359 6 364 147
rect 99 3 364 6
<< metal2 >>
rect 88 119 168 122
rect 88 113 91 119
rect 49 110 91 113
rect 164 112 167 119
rect 188 117 247 120
rect 121 109 142 112
rect 168 109 194 112
rect 198 109 199 112
rect 244 111 247 117
rect 268 112 287 115
rect 244 108 251 111
rect 268 107 271 112
rect 291 113 330 114
rect 291 111 326 113
rect 64 99 76 102
rect 73 35 76 99
rect 136 99 218 102
rect 281 102 340 105
rect 251 97 254 100
rect 251 94 309 97
rect 240 75 244 93
rect 121 71 244 75
rect 121 45 125 71
rect 240 70 244 71
rect 255 56 313 59
rect 140 51 222 54
rect 255 53 258 56
rect 285 48 344 51
rect 125 41 146 44
rect 172 41 198 44
rect 202 41 203 44
rect 248 42 255 45
rect 168 35 171 41
rect 73 32 171 35
rect 248 36 251 42
rect 295 40 330 42
rect 295 39 334 40
rect 192 33 251 36
<< ntransistor >>
rect 40 87 42 90
rect 112 86 114 89
rect 151 86 153 92
rect 172 86 174 92
rect 205 86 207 92
rect 226 86 228 92
rect 261 86 263 92
rect 282 86 284 92
rect 315 86 317 92
rect 336 86 338 92
rect 116 64 118 67
rect 155 61 157 67
rect 176 61 178 67
rect 209 61 211 67
rect 230 61 232 67
rect 265 61 267 67
rect 286 61 288 67
rect 319 61 321 67
rect 340 61 342 67
<< ptransistor >>
rect 40 123 42 129
rect 112 123 114 129
rect 151 123 153 129
rect 172 123 174 129
rect 205 123 207 129
rect 226 123 228 129
rect 261 123 263 129
rect 282 123 284 129
rect 315 123 317 129
rect 336 123 338 129
rect 116 24 118 30
rect 155 24 157 30
rect 176 24 178 30
rect 209 24 211 30
rect 230 24 232 30
rect 265 24 267 30
rect 286 24 288 30
rect 319 24 321 30
rect 340 24 342 30
<< polycontact >>
rect 38 108 42 112
rect 110 107 114 111
rect 148 107 152 111
rect 169 107 173 111
rect 202 107 206 111
rect 223 107 227 111
rect 258 107 262 111
rect 279 107 283 111
rect 312 107 316 111
rect 333 107 337 111
rect 114 42 118 46
rect 152 42 156 46
rect 173 42 177 46
rect 206 42 210 46
rect 227 42 231 46
rect 262 42 266 46
rect 283 42 287 46
rect 316 42 320 46
rect 337 42 341 46
<< ndcontact >>
rect 25 87 29 91
rect 59 87 63 91
rect 97 86 101 90
rect 131 86 135 90
rect 143 87 147 91
rect 177 87 181 91
rect 197 87 201 91
rect 231 87 235 91
rect 253 87 257 91
rect 287 87 291 91
rect 307 87 311 91
rect 341 87 345 91
rect 101 63 105 67
rect 135 63 139 67
rect 147 62 151 66
rect 181 62 185 66
rect 201 62 205 66
rect 235 62 239 66
rect 257 62 261 66
rect 291 62 295 66
rect 311 62 315 66
rect 345 62 349 66
<< pdcontact >>
rect 14 124 18 128
rect 58 124 64 130
rect 97 124 101 128
rect 130 124 134 128
rect 143 124 147 128
rect 160 124 164 128
rect 177 124 181 128
rect 197 124 201 128
rect 214 124 218 128
rect 231 124 235 128
rect 253 124 257 128
rect 270 124 274 128
rect 287 124 291 128
rect 307 124 311 128
rect 324 124 328 128
rect 341 124 345 128
rect 101 25 105 29
rect 134 25 138 29
rect 147 25 151 29
rect 164 25 168 29
rect 181 25 185 29
rect 201 25 205 29
rect 218 25 222 29
rect 235 25 239 29
rect 257 25 261 29
rect 274 25 278 29
rect 291 25 295 29
rect 311 25 315 29
rect 328 25 332 29
rect 345 25 349 29
<< m2contact >>
rect 45 109 49 113
rect 117 108 121 112
rect 60 99 64 103
rect 142 108 146 112
rect 164 108 168 112
rect 184 116 188 120
rect 194 108 198 112
rect 132 98 136 102
rect 218 99 222 103
rect 251 108 255 112
rect 287 111 291 115
rect 250 100 254 104
rect 267 103 271 107
rect 277 101 281 105
rect 240 93 244 97
rect 326 109 330 113
rect 340 102 344 106
rect 309 94 313 98
rect 136 51 140 55
rect 121 41 125 45
rect 222 50 226 54
rect 254 49 258 53
rect 146 41 150 45
rect 168 41 172 45
rect 198 41 202 45
rect 281 48 285 52
rect 255 41 259 45
rect 313 55 317 59
rect 344 47 348 51
rect 291 38 295 42
rect 330 40 334 44
rect 188 33 192 37
<< nsubstratencontact >>
rect 170 138 174 142
rect 224 138 228 142
rect 280 138 284 142
rect 334 138 338 142
rect 174 11 178 15
rect 228 11 232 15
rect 284 11 288 15
rect 338 11 342 15
<< labels >>
rlabel metal1 330 5 330 5 1 vdd
rlabel ndiffusion 330 64 330 64 1 n10
rlabel m2contact 61 101 61 101 1 en_bar_D3
rlabel metal1 132 108 132 108 1 D_bar_D3
rlabel polycontact 150 109 150 109 1 D_D3
rlabel polycontact 171 109 171 109 1 en_D3
rlabel ndiffusion 160 89 160 89 1 n1_D3
rlabel metal1 179 106 179 106 1 out_n1_D3
rlabel ndiffusion 216 89 216 89 1 n2_D3
rlabel metal1 234 102 234 102 1 out_n2_D3
rlabel ndiffusion 272 89 272 89 1 n3_D3
rlabel ndiffusion 326 89 326 89 1 n4_D3
rlabel m2contact 343 105 343 105 1 q_l1_bar_D3
rlabel m2contact 347 48 347 48 1 q_bar_D3
rlabel ndiffusion 276 64 276 64 1 n9_D3
rlabel metal1 238 51 238 51 1 out_n8_D3
rlabel m2contact 293 40 293 40 1 q_D3
rlabel ndiffusion 220 64 220 64 1 n8_D3
rlabel metal1 183 47 183 47 1 out_n7_D3
rlabel ndiffusion 164 64 164 64 1 n7_D3
rlabel polycontact 154 44 154 44 1 q_l1_D3
rlabel metal1 136 48 136 48 1 n6_D3
rlabel metal1 171 79 171 79 1 vss
<< end >>
