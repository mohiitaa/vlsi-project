magic
tech scmos
timestamp 1523162757
<< pwell >>
rect 110 457 128 461
rect 108 453 128 457
rect 108 417 156 453
rect 195 417 243 453
rect 288 417 336 453
rect 528 419 576 455
rect 621 419 669 455
rect 708 419 756 455
rect 37 294 180 330
rect 192 294 310 330
rect 366 296 509 332
rect 521 296 639 332
rect 693 299 836 335
rect 1563 358 1599 444
rect 848 299 966 335
rect 123 268 171 294
rect 452 270 500 296
rect 779 273 827 299
rect 1537 310 1599 358
rect 1687 362 1723 480
rect 1687 357 1711 362
rect 1689 350 1711 357
rect 1689 341 1723 350
rect 1563 301 1599 310
rect 1687 293 1749 341
rect 1370 245 1410 270
rect 1370 234 1411 245
rect 36 148 179 184
rect 191 148 309 184
rect 365 150 508 186
rect 520 150 638 186
rect 692 153 835 189
rect 1371 209 1411 234
rect 847 153 965 189
rect 122 122 170 148
rect 451 124 499 150
rect 778 127 826 153
rect 1563 171 1599 289
rect 1687 207 1723 293
rect 1370 94 1411 130
rect 323 0 371 36
rect 416 0 464 36
rect 503 0 551 36
rect 1565 -2 1601 84
rect 121 -49 139 -45
rect 119 -53 139 -49
rect 1539 -50 1601 -2
rect 1689 2 1725 120
rect 1689 -3 1713 2
rect 1691 -10 1713 -3
rect 1691 -19 1725 -10
rect 119 -89 167 -53
rect 206 -89 254 -53
rect 299 -89 347 -53
rect 539 -87 587 -51
rect 632 -87 680 -51
rect 719 -87 767 -51
rect 1565 -59 1601 -50
rect 1689 -67 1751 -19
rect 48 -212 191 -176
rect 203 -212 321 -176
rect 377 -210 520 -174
rect 532 -210 650 -174
rect 704 -207 847 -171
rect 859 -207 977 -171
rect 1565 -189 1601 -71
rect 1689 -153 1725 -67
rect 134 -238 182 -212
rect 463 -236 511 -210
rect 790 -233 838 -207
rect 1402 -264 1442 -228
rect 47 -358 190 -322
rect 202 -358 320 -322
rect 376 -356 519 -320
rect 531 -356 649 -320
rect 703 -353 846 -317
rect 858 -353 976 -317
rect 133 -384 181 -358
rect 462 -382 510 -356
rect 789 -379 837 -353
rect 1681 -354 1717 -236
rect 1404 -397 1444 -365
rect 1404 -407 1445 -397
rect 1404 -409 1446 -407
rect 334 -506 382 -470
rect 427 -506 475 -470
rect 1406 -443 1446 -409
rect 514 -506 562 -470
rect 1681 -375 1717 -366
rect 1681 -418 1743 -375
rect 1681 -509 1742 -418
rect 1706 -527 1742 -509
<< nwell >>
rect 1643 479 1687 480
rect 108 374 156 417
rect 195 374 243 417
rect 288 374 336 417
rect 528 382 576 419
rect 621 382 669 419
rect 528 379 669 382
rect 524 376 669 379
rect 1005 421 1184 447
rect 1197 421 1238 447
rect 1253 421 1294 447
rect 1307 421 1348 447
rect 1636 444 1687 479
rect 708 388 756 419
rect 708 379 769 388
rect 708 376 836 379
rect 37 330 180 374
rect 192 373 336 374
rect 192 330 310 373
rect 366 332 509 376
rect 521 362 836 376
rect 521 332 639 362
rect 693 335 836 362
rect 848 335 966 379
rect 1517 358 1530 362
rect 1101 316 1188 342
rect 1201 316 1242 342
rect 1257 316 1298 342
rect 1311 316 1352 342
rect 123 261 171 268
rect 452 263 500 270
rect 1005 276 1184 302
rect 1197 276 1238 302
rect 1253 276 1294 302
rect 1307 276 1348 302
rect 779 266 827 273
rect 119 248 171 261
rect 448 250 500 263
rect 775 253 827 266
rect 123 232 171 248
rect 452 234 500 250
rect 779 240 827 253
rect 1370 270 1410 314
rect 1494 310 1537 358
rect 1599 357 1687 444
rect 1599 341 1689 357
rect 1599 301 1687 341
rect 1639 289 1687 301
rect 1749 293 1793 341
rect 112 228 178 232
rect 442 230 508 234
rect 750 233 861 240
rect 36 184 179 228
rect 191 184 309 228
rect 365 186 508 230
rect 520 186 638 230
rect 692 224 965 233
rect 692 189 835 224
rect 847 189 965 224
rect 1101 171 1188 197
rect 1201 171 1242 197
rect 1257 171 1298 197
rect 1311 174 1352 197
rect 1371 174 1411 209
rect 1340 171 1352 174
rect 122 115 170 122
rect 451 117 499 124
rect 1004 134 1183 160
rect 1196 134 1237 160
rect 1252 134 1293 160
rect 1306 134 1347 160
rect 778 120 826 127
rect 118 102 170 115
rect 447 104 499 117
rect 774 107 826 120
rect 122 78 170 102
rect 451 94 499 104
rect 325 80 557 94
rect 778 83 826 107
rect 1370 130 1411 174
rect 1599 207 1687 289
rect 1756 289 1769 293
rect 1599 173 1648 207
rect 1599 171 1643 173
rect 1645 119 1689 120
rect 1638 84 1689 119
rect 323 77 557 80
rect 323 36 371 77
rect 416 36 464 77
rect 503 36 551 77
rect 1100 29 1187 55
rect 1200 29 1241 55
rect 1256 29 1297 55
rect 1310 29 1351 55
rect 1519 -2 1532 2
rect 1496 -50 1539 -2
rect 1601 -3 1689 84
rect 1601 -19 1691 -3
rect 119 -132 167 -89
rect 206 -132 254 -89
rect 299 -132 347 -89
rect 539 -124 587 -87
rect 632 -124 680 -87
rect 539 -127 680 -124
rect 535 -130 680 -127
rect 1601 -59 1689 -19
rect 719 -118 767 -87
rect 1026 -90 1205 -64
rect 1218 -90 1259 -64
rect 1274 -90 1315 -64
rect 1328 -90 1369 -64
rect 1641 -71 1689 -59
rect 1751 -67 1795 -19
rect 719 -127 780 -118
rect 719 -130 847 -127
rect 48 -176 191 -132
rect 203 -133 347 -132
rect 203 -176 321 -133
rect 377 -174 520 -130
rect 532 -144 847 -130
rect 532 -174 650 -144
rect 704 -171 847 -144
rect 859 -171 977 -127
rect 1122 -195 1209 -169
rect 1222 -195 1263 -169
rect 1278 -195 1319 -169
rect 1332 -195 1373 -169
rect 1601 -153 1689 -71
rect 1758 -71 1771 -67
rect 1601 -187 1650 -153
rect 1601 -189 1645 -187
rect 134 -245 182 -238
rect 463 -243 511 -236
rect 790 -240 838 -233
rect 1024 -235 1203 -209
rect 1216 -235 1257 -209
rect 1272 -235 1313 -209
rect 1326 -235 1367 -209
rect 130 -258 182 -245
rect 459 -256 511 -243
rect 786 -253 838 -240
rect 134 -274 182 -258
rect 463 -272 511 -256
rect 790 -266 838 -253
rect 123 -278 189 -274
rect 453 -276 519 -272
rect 761 -273 872 -266
rect 47 -322 190 -278
rect 202 -322 320 -278
rect 376 -320 519 -276
rect 531 -320 649 -276
rect 703 -282 976 -273
rect 703 -317 846 -282
rect 858 -317 976 -282
rect 1402 -305 1442 -264
rect 1401 -308 1442 -305
rect 1120 -340 1207 -314
rect 1220 -340 1261 -314
rect 1276 -340 1317 -314
rect 1330 -340 1371 -314
rect 1401 -321 1441 -308
rect 133 -391 181 -384
rect 462 -389 510 -382
rect 1025 -377 1204 -351
rect 1217 -377 1258 -351
rect 1273 -377 1314 -351
rect 1327 -377 1368 -351
rect 1404 -365 1444 -321
rect 1637 -354 1681 -236
rect 789 -386 837 -379
rect 129 -404 181 -391
rect 458 -402 510 -389
rect 785 -399 837 -386
rect 133 -428 181 -404
rect 462 -412 510 -402
rect 336 -426 568 -412
rect 789 -423 837 -399
rect 334 -429 568 -426
rect 334 -470 382 -429
rect 427 -470 475 -429
rect 514 -470 562 -429
rect 1121 -482 1208 -456
rect 1221 -482 1262 -456
rect 1277 -482 1318 -456
rect 1331 -482 1372 -456
rect 1406 -487 1446 -443
rect 1637 -509 1681 -366
rect 1743 -418 1787 -375
rect 1742 -423 1787 -418
rect 1742 -527 1786 -423
<< polysilicon >>
rect 1692 469 1698 470
rect 1692 467 1693 469
rect 1666 465 1671 467
rect 1681 465 1693 467
rect 1697 466 1698 469
rect 1697 465 1701 466
rect 1692 464 1701 465
rect 1710 464 1715 466
rect 1660 460 1666 461
rect 1660 456 1661 460
rect 1665 457 1666 460
rect 1684 457 1701 459
rect 1710 457 1715 459
rect 1665 456 1671 457
rect 1660 455 1671 456
rect 1681 455 1687 457
rect 121 436 123 441
rect 128 436 130 441
rect 141 434 143 438
rect 208 436 210 441
rect 215 436 217 441
rect 228 434 230 438
rect 301 436 303 441
rect 308 436 310 441
rect 321 434 323 438
rect 541 436 543 440
rect 554 438 556 443
rect 561 438 563 443
rect 634 436 636 440
rect 647 438 649 443
rect 654 438 656 443
rect 721 436 723 440
rect 734 438 736 443
rect 741 438 743 443
rect 1042 434 1044 436
rect 1114 434 1116 440
rect 1153 434 1155 440
rect 1174 434 1176 440
rect 1207 434 1209 440
rect 1228 434 1230 440
rect 1263 434 1265 440
rect 1284 434 1286 440
rect 1317 434 1319 440
rect 1338 434 1340 440
rect 1684 450 1690 451
rect 1684 447 1685 450
rect 1664 445 1669 447
rect 1681 446 1685 447
rect 1689 447 1690 450
rect 1689 446 1698 447
rect 1681 445 1698 446
rect 1704 445 1708 447
rect 1578 436 1582 438
rect 1588 437 1605 438
rect 1588 436 1597 437
rect 1596 433 1597 436
rect 1601 436 1605 437
rect 1617 436 1622 438
rect 1601 433 1602 436
rect 1596 432 1602 433
rect 121 412 123 425
rect 128 420 130 425
rect 141 420 143 425
rect 127 419 133 420
rect 127 415 128 419
rect 132 415 133 419
rect 127 414 133 415
rect 137 419 143 420
rect 137 415 138 419
rect 142 415 143 419
rect 137 414 143 415
rect 117 411 123 412
rect 117 407 118 411
rect 122 407 123 411
rect 117 406 123 407
rect 121 403 123 406
rect 131 403 133 414
rect 141 410 143 414
rect 208 412 210 425
rect 215 420 217 425
rect 228 420 230 425
rect 214 419 220 420
rect 214 415 215 419
rect 219 415 220 419
rect 214 414 220 415
rect 224 419 230 420
rect 224 415 225 419
rect 229 415 230 419
rect 224 414 230 415
rect 204 411 210 412
rect 204 407 205 411
rect 209 407 210 411
rect 204 406 210 407
rect 208 403 210 406
rect 218 403 220 414
rect 228 410 230 414
rect 301 412 303 425
rect 308 420 310 425
rect 321 420 323 425
rect 307 419 313 420
rect 307 415 308 419
rect 312 415 313 419
rect 307 414 313 415
rect 317 419 323 420
rect 317 415 318 419
rect 322 415 323 419
rect 317 414 323 415
rect 297 411 303 412
rect 121 385 123 390
rect 131 385 133 390
rect 141 388 143 392
rect 297 407 298 411
rect 302 407 303 411
rect 297 406 303 407
rect 301 403 303 406
rect 311 403 313 414
rect 321 410 323 414
rect 541 422 543 427
rect 554 422 556 427
rect 541 421 547 422
rect 541 417 542 421
rect 546 417 547 421
rect 541 416 547 417
rect 551 421 557 422
rect 551 417 552 421
rect 556 417 557 421
rect 551 416 557 417
rect 541 412 543 416
rect 208 385 210 390
rect 218 385 220 390
rect 228 388 230 392
rect 551 405 553 416
rect 561 414 563 427
rect 634 422 636 427
rect 647 422 649 427
rect 634 421 640 422
rect 634 417 635 421
rect 639 417 640 421
rect 634 416 640 417
rect 644 421 650 422
rect 644 417 645 421
rect 649 417 650 421
rect 644 416 650 417
rect 561 413 567 414
rect 561 409 562 413
rect 566 409 567 413
rect 634 412 636 416
rect 561 408 567 409
rect 561 405 563 408
rect 301 385 303 390
rect 311 385 313 390
rect 321 388 323 392
rect 541 390 543 394
rect 644 405 646 416
rect 654 414 656 427
rect 721 422 723 427
rect 734 422 736 427
rect 721 421 727 422
rect 721 417 722 421
rect 726 417 727 421
rect 721 416 727 417
rect 731 421 737 422
rect 731 417 732 421
rect 736 417 737 421
rect 731 416 737 417
rect 654 413 660 414
rect 654 409 655 413
rect 659 409 660 413
rect 721 412 723 416
rect 654 408 660 409
rect 654 405 656 408
rect 551 387 553 392
rect 561 387 563 392
rect 634 390 636 394
rect 731 405 733 416
rect 741 414 743 427
rect 1042 417 1044 428
rect 741 413 747 414
rect 1114 416 1116 428
rect 1153 416 1155 428
rect 1174 416 1176 428
rect 1207 416 1209 428
rect 1228 416 1230 428
rect 1263 416 1265 428
rect 1284 416 1286 428
rect 1317 416 1319 428
rect 1338 416 1340 428
rect 1599 426 1605 428
rect 1615 427 1626 428
rect 1615 426 1621 427
rect 1571 424 1576 426
rect 1585 424 1602 426
rect 1620 423 1621 426
rect 1625 423 1626 427
rect 1620 422 1626 423
rect 1571 417 1576 419
rect 1585 418 1594 419
rect 1585 417 1589 418
rect 741 409 742 413
rect 746 409 747 413
rect 741 408 747 409
rect 741 405 743 408
rect 644 387 646 392
rect 654 387 656 392
rect 721 390 723 394
rect 1042 395 1044 413
rect 1154 412 1155 416
rect 1175 412 1176 416
rect 1208 412 1209 416
rect 1229 412 1230 416
rect 1264 412 1265 416
rect 1285 412 1286 416
rect 1318 412 1319 416
rect 1339 412 1340 416
rect 731 387 733 392
rect 741 387 743 392
rect 1042 389 1044 392
rect 1114 394 1116 412
rect 1153 397 1155 412
rect 1174 397 1176 412
rect 1207 397 1209 412
rect 1228 397 1230 412
rect 1263 397 1265 412
rect 1284 397 1286 412
rect 1317 397 1319 412
rect 1338 397 1340 412
rect 1588 414 1589 417
rect 1593 416 1605 418
rect 1615 416 1620 418
rect 1593 414 1594 416
rect 1588 413 1594 414
rect 1649 419 1653 421
rect 1680 420 1689 421
rect 1680 419 1684 420
rect 1683 416 1684 419
rect 1688 418 1698 420
rect 1710 418 1715 420
rect 1688 416 1689 418
rect 1683 415 1689 416
rect 1693 411 1698 413
rect 1710 411 1715 413
rect 1658 409 1662 411
rect 1680 410 1695 411
rect 1680 409 1684 410
rect 1683 406 1684 409
rect 1688 409 1695 410
rect 1688 406 1689 409
rect 1683 405 1689 406
rect 1693 401 1698 403
rect 1707 401 1717 403
rect 1658 399 1662 401
rect 1680 399 1685 401
rect 1683 393 1685 399
rect 1683 391 1698 393
rect 1707 391 1711 393
rect 1114 388 1116 391
rect 1153 388 1155 391
rect 1174 388 1176 391
rect 1207 388 1209 391
rect 1228 388 1230 391
rect 1263 388 1265 391
rect 1284 388 1286 391
rect 1317 388 1319 391
rect 1338 388 1340 391
rect 1689 389 1695 391
rect 1689 385 1690 389
rect 1694 385 1695 389
rect 1649 383 1653 385
rect 1680 383 1685 385
rect 1689 384 1695 385
rect 1683 377 1685 383
rect 1715 380 1717 401
rect 1705 378 1717 380
rect 1705 377 1707 378
rect 1683 375 1693 377
rect 1702 375 1707 377
rect 129 364 131 368
rect 53 356 59 357
rect 43 348 45 353
rect 53 352 54 356
rect 58 352 59 356
rect 53 351 59 352
rect 53 346 55 351
rect 63 346 65 351
rect 114 348 120 349
rect 114 344 115 348
rect 119 344 120 348
rect 114 343 120 344
rect 43 333 45 336
rect 53 333 55 336
rect 43 332 49 333
rect 43 328 44 332
rect 48 328 49 332
rect 53 330 57 333
rect 43 327 49 328
rect 43 319 45 327
rect 55 316 57 330
rect 63 325 65 336
rect 118 334 120 343
rect 165 364 167 368
rect 213 364 215 368
rect 145 355 147 359
rect 155 355 157 359
rect 198 348 204 349
rect 198 344 199 348
rect 203 344 204 348
rect 198 343 204 344
rect 129 334 131 337
rect 145 334 147 337
rect 155 334 157 337
rect 165 334 167 337
rect 118 332 131 334
rect 137 332 147 334
rect 151 333 157 334
rect 62 324 68 325
rect 121 324 123 332
rect 137 328 139 332
rect 151 329 152 333
rect 156 329 157 333
rect 151 328 157 329
rect 161 333 167 334
rect 161 329 162 333
rect 166 329 167 333
rect 202 334 204 343
rect 249 364 251 368
rect 229 355 231 359
rect 239 355 241 359
rect 458 366 460 370
rect 382 358 388 359
rect 285 356 291 357
rect 275 348 277 353
rect 285 352 286 356
rect 290 352 291 356
rect 285 351 291 352
rect 213 334 215 337
rect 229 334 231 337
rect 239 334 241 337
rect 249 334 251 337
rect 285 346 287 351
rect 295 346 297 351
rect 372 350 374 355
rect 382 354 383 358
rect 387 354 388 358
rect 382 353 388 354
rect 382 348 384 353
rect 392 348 394 353
rect 443 350 449 351
rect 443 346 444 350
rect 448 346 449 350
rect 443 345 449 346
rect 202 332 215 334
rect 221 332 231 334
rect 235 333 241 334
rect 161 328 167 329
rect 130 327 139 328
rect 62 320 63 324
rect 67 320 68 324
rect 62 319 68 320
rect 62 316 64 319
rect 43 309 45 313
rect 130 323 131 327
rect 135 323 139 327
rect 155 324 157 328
rect 130 322 139 323
rect 137 319 139 322
rect 147 319 149 324
rect 155 322 159 324
rect 157 319 159 322
rect 164 319 166 328
rect 205 324 207 332
rect 221 328 223 332
rect 235 329 236 333
rect 240 329 241 333
rect 235 328 241 329
rect 245 333 251 334
rect 245 329 246 333
rect 250 329 251 333
rect 245 328 251 329
rect 275 333 277 336
rect 285 333 287 336
rect 275 332 281 333
rect 275 328 276 332
rect 280 328 281 332
rect 285 330 289 333
rect 214 327 223 328
rect 121 312 123 315
rect 121 310 126 312
rect 55 302 57 307
rect 62 302 64 307
rect 124 302 126 310
rect 137 306 139 310
rect 147 302 149 310
rect 214 323 215 327
rect 219 323 223 327
rect 239 324 241 328
rect 214 322 223 323
rect 221 319 223 322
rect 231 319 233 324
rect 239 322 243 324
rect 241 319 243 322
rect 248 319 250 328
rect 275 327 281 328
rect 275 319 277 327
rect 205 312 207 315
rect 205 310 210 312
rect 157 302 159 307
rect 164 302 166 307
rect 124 300 149 302
rect 208 302 210 310
rect 221 306 223 310
rect 231 302 233 310
rect 287 316 289 330
rect 295 325 297 336
rect 372 335 374 338
rect 382 335 384 338
rect 372 334 378 335
rect 372 330 373 334
rect 377 330 378 334
rect 382 332 386 335
rect 372 329 378 330
rect 294 324 300 325
rect 294 320 295 324
rect 299 320 300 324
rect 372 321 374 329
rect 294 319 300 320
rect 294 316 296 319
rect 275 309 277 313
rect 384 318 386 332
rect 392 327 394 338
rect 447 336 449 345
rect 494 366 496 370
rect 542 366 544 370
rect 474 357 476 361
rect 484 357 486 361
rect 527 350 533 351
rect 527 346 528 350
rect 532 346 533 350
rect 527 345 533 346
rect 458 336 460 339
rect 474 336 476 339
rect 484 336 486 339
rect 494 336 496 339
rect 447 334 460 336
rect 466 334 476 336
rect 480 335 486 336
rect 391 326 397 327
rect 450 326 452 334
rect 466 330 468 334
rect 480 331 481 335
rect 485 331 486 335
rect 480 330 486 331
rect 490 335 496 336
rect 490 331 491 335
rect 495 331 496 335
rect 531 336 533 345
rect 578 366 580 370
rect 558 357 560 361
rect 568 357 570 361
rect 785 369 787 373
rect 709 361 715 362
rect 614 358 620 359
rect 604 350 606 355
rect 614 354 615 358
rect 619 354 620 358
rect 614 353 620 354
rect 699 353 701 358
rect 709 357 710 361
rect 714 357 715 361
rect 709 356 715 357
rect 542 336 544 339
rect 558 336 560 339
rect 568 336 570 339
rect 578 336 580 339
rect 614 348 616 353
rect 624 348 626 353
rect 709 351 711 356
rect 719 351 721 356
rect 770 353 776 354
rect 770 349 771 353
rect 775 349 776 353
rect 770 348 776 349
rect 699 338 701 341
rect 709 338 711 341
rect 531 334 544 336
rect 550 334 560 336
rect 564 335 570 336
rect 490 330 496 331
rect 459 329 468 330
rect 391 322 392 326
rect 396 322 397 326
rect 391 321 397 322
rect 391 318 393 321
rect 372 311 374 315
rect 459 325 460 329
rect 464 325 468 329
rect 484 326 486 330
rect 459 324 468 325
rect 466 321 468 324
rect 476 321 478 326
rect 484 324 488 326
rect 486 321 488 324
rect 493 321 495 330
rect 534 326 536 334
rect 550 330 552 334
rect 564 331 565 335
rect 569 331 570 335
rect 564 330 570 331
rect 574 335 580 336
rect 574 331 575 335
rect 579 331 580 335
rect 574 330 580 331
rect 604 335 606 338
rect 614 335 616 338
rect 604 334 610 335
rect 604 330 605 334
rect 609 330 610 334
rect 614 332 618 335
rect 543 329 552 330
rect 450 314 452 317
rect 450 312 455 314
rect 241 302 243 307
rect 248 302 250 307
rect 208 300 233 302
rect 287 302 289 307
rect 294 302 296 307
rect 384 304 386 309
rect 391 304 393 309
rect 453 304 455 312
rect 466 308 468 312
rect 476 304 478 312
rect 543 325 544 329
rect 548 325 552 329
rect 568 326 570 330
rect 543 324 552 325
rect 550 321 552 324
rect 560 321 562 326
rect 568 324 572 326
rect 570 321 572 324
rect 577 321 579 330
rect 604 329 610 330
rect 604 321 606 329
rect 534 314 536 317
rect 534 312 539 314
rect 486 304 488 309
rect 493 304 495 309
rect 453 302 478 304
rect 537 304 539 312
rect 550 308 552 312
rect 560 304 562 312
rect 616 318 618 332
rect 624 327 626 338
rect 699 337 705 338
rect 699 333 700 337
rect 704 333 705 337
rect 709 335 713 338
rect 699 332 705 333
rect 623 326 629 327
rect 623 322 624 326
rect 628 322 629 326
rect 699 324 701 332
rect 623 321 629 322
rect 623 318 625 321
rect 711 321 713 335
rect 719 330 721 341
rect 774 339 776 348
rect 821 369 823 373
rect 869 369 871 373
rect 801 360 803 364
rect 811 360 813 364
rect 854 353 860 354
rect 854 349 855 353
rect 859 349 860 353
rect 854 348 860 349
rect 785 339 787 342
rect 801 339 803 342
rect 811 339 813 342
rect 821 339 823 342
rect 774 337 787 339
rect 793 337 803 339
rect 807 338 813 339
rect 718 329 724 330
rect 777 329 779 337
rect 793 333 795 337
rect 807 334 808 338
rect 812 334 813 338
rect 807 333 813 334
rect 817 338 823 339
rect 817 334 818 338
rect 822 334 823 338
rect 858 339 860 348
rect 905 369 907 373
rect 1118 372 1120 375
rect 1157 372 1159 375
rect 1178 372 1180 375
rect 1211 372 1213 375
rect 1232 372 1234 375
rect 1267 372 1269 375
rect 1288 372 1290 375
rect 1321 372 1323 375
rect 1342 372 1344 375
rect 1683 374 1685 375
rect 1668 373 1685 374
rect 885 360 887 364
rect 895 360 897 364
rect 941 361 947 362
rect 931 353 933 358
rect 941 357 942 361
rect 946 357 947 361
rect 941 356 947 357
rect 869 339 871 342
rect 885 339 887 342
rect 895 339 897 342
rect 905 339 907 342
rect 941 351 943 356
rect 951 351 953 356
rect 1118 351 1120 369
rect 1668 369 1669 373
rect 1673 372 1685 373
rect 1673 369 1674 372
rect 1668 368 1674 369
rect 1157 351 1159 366
rect 1178 351 1180 366
rect 1211 351 1213 366
rect 1232 351 1234 366
rect 1267 351 1269 366
rect 1288 351 1290 366
rect 1321 351 1323 366
rect 1342 351 1344 366
rect 1612 366 1618 367
rect 1612 363 1613 366
rect 1601 362 1613 363
rect 1617 362 1618 366
rect 1601 361 1618 362
rect 1601 360 1603 361
rect 1579 358 1584 360
rect 1593 358 1603 360
rect 1579 357 1581 358
rect 1569 355 1581 357
rect 1158 347 1159 351
rect 1179 347 1180 351
rect 1212 347 1213 351
rect 1233 347 1234 351
rect 1268 347 1269 351
rect 1289 347 1290 351
rect 1322 347 1323 351
rect 1343 347 1344 351
rect 858 337 871 339
rect 877 337 887 339
rect 891 338 897 339
rect 817 333 823 334
rect 786 332 795 333
rect 718 325 719 329
rect 723 325 724 329
rect 718 324 724 325
rect 718 321 720 324
rect 604 311 606 315
rect 699 314 701 318
rect 786 328 787 332
rect 791 328 795 332
rect 811 329 813 333
rect 786 327 795 328
rect 793 324 795 327
rect 803 324 805 329
rect 811 327 815 329
rect 813 324 815 327
rect 820 324 822 333
rect 861 329 863 337
rect 877 333 879 337
rect 891 334 892 338
rect 896 334 897 338
rect 891 333 897 334
rect 901 338 907 339
rect 901 334 902 338
rect 906 334 907 338
rect 901 333 907 334
rect 931 338 933 341
rect 941 338 943 341
rect 931 337 937 338
rect 931 333 932 337
rect 936 333 937 337
rect 941 335 945 338
rect 870 332 879 333
rect 777 317 779 320
rect 777 315 782 317
rect 570 304 572 309
rect 577 304 579 309
rect 537 302 562 304
rect 616 304 618 309
rect 623 304 625 309
rect 711 307 713 312
rect 718 307 720 312
rect 780 307 782 315
rect 793 311 795 315
rect 803 307 805 315
rect 870 328 871 332
rect 875 328 879 332
rect 895 329 897 333
rect 870 327 879 328
rect 877 324 879 327
rect 887 324 889 329
rect 895 327 899 329
rect 897 324 899 327
rect 904 324 906 333
rect 931 332 937 333
rect 931 324 933 332
rect 861 317 863 320
rect 861 315 866 317
rect 813 307 815 312
rect 820 307 822 312
rect 780 305 805 307
rect 864 307 866 315
rect 877 311 879 315
rect 887 307 889 315
rect 943 321 945 335
rect 951 330 953 341
rect 1118 335 1120 347
rect 1157 335 1159 347
rect 1178 335 1180 347
rect 1211 335 1213 347
rect 1232 335 1234 347
rect 1267 335 1269 347
rect 1288 335 1290 347
rect 1321 335 1323 347
rect 1342 335 1344 347
rect 1534 348 1540 349
rect 1534 345 1535 348
rect 1499 343 1503 345
rect 1521 344 1535 345
rect 1539 345 1540 348
rect 1539 344 1548 345
rect 1521 343 1548 344
rect 1554 343 1558 345
rect 1526 338 1532 339
rect 1499 336 1503 338
rect 1521 336 1527 338
rect 950 329 956 330
rect 1526 334 1527 336
rect 1531 335 1532 338
rect 1531 334 1535 335
rect 1526 333 1535 334
rect 1539 333 1548 335
rect 1554 333 1558 335
rect 950 325 951 329
rect 955 325 956 329
rect 950 324 956 325
rect 950 321 952 324
rect 1118 323 1120 329
rect 1157 323 1159 329
rect 1178 323 1180 329
rect 1211 323 1213 329
rect 1232 323 1234 329
rect 1267 323 1269 329
rect 1288 323 1290 329
rect 1321 323 1323 329
rect 1342 323 1344 329
rect 1533 328 1539 329
rect 1533 325 1534 328
rect 1508 323 1512 325
rect 1524 324 1534 325
rect 1538 325 1539 328
rect 1538 324 1548 325
rect 1524 323 1548 324
rect 1554 323 1558 325
rect 931 314 933 318
rect 1569 334 1571 355
rect 1601 352 1603 358
rect 1591 350 1597 351
rect 1601 350 1606 352
rect 1633 350 1637 352
rect 1591 346 1592 350
rect 1596 346 1597 350
rect 1591 344 1597 346
rect 1575 342 1579 344
rect 1588 342 1603 344
rect 1601 336 1603 342
rect 1601 334 1606 336
rect 1624 334 1628 336
rect 1649 335 1653 337
rect 1680 336 1689 337
rect 1680 335 1684 336
rect 1569 332 1579 334
rect 1588 332 1593 334
rect 1597 329 1603 330
rect 1597 326 1598 329
rect 1591 325 1598 326
rect 1602 326 1603 329
rect 1683 332 1684 335
rect 1688 334 1698 336
rect 1710 334 1715 336
rect 1688 332 1689 334
rect 1683 331 1689 332
rect 1693 327 1698 329
rect 1710 327 1715 329
rect 1602 325 1606 326
rect 1591 324 1606 325
rect 1624 324 1628 326
rect 1658 325 1662 327
rect 1680 326 1695 327
rect 1680 325 1684 326
rect 1571 322 1576 324
rect 1588 322 1593 324
rect 1597 319 1603 320
rect 1597 317 1598 319
rect 1571 315 1576 317
rect 1588 315 1598 317
rect 1602 316 1603 319
rect 1683 322 1684 325
rect 1688 325 1695 326
rect 1688 322 1689 325
rect 1683 321 1689 322
rect 1693 317 1698 319
rect 1707 317 1717 319
rect 1602 315 1606 316
rect 1597 314 1606 315
rect 1633 314 1637 316
rect 1658 315 1662 317
rect 1680 315 1685 317
rect 897 307 899 312
rect 904 307 906 312
rect 864 305 889 307
rect 943 307 945 312
rect 950 307 952 312
rect 1395 304 1397 308
rect 1683 309 1685 315
rect 1683 307 1698 309
rect 1707 307 1711 309
rect 136 285 138 289
rect 146 285 148 289
rect 156 285 158 289
rect 465 287 467 291
rect 475 287 477 291
rect 485 287 487 291
rect 792 290 794 294
rect 802 290 804 294
rect 812 290 814 294
rect 1042 289 1044 291
rect 136 271 138 279
rect 132 270 138 271
rect 146 270 148 279
rect 156 270 158 279
rect 465 273 467 281
rect 132 266 133 270
rect 137 266 138 270
rect 152 269 158 270
rect 132 265 138 266
rect 136 252 138 265
rect 146 263 148 266
rect 152 265 153 269
rect 157 265 158 269
rect 461 272 467 273
rect 475 272 477 281
rect 485 272 487 281
rect 792 276 794 284
rect 461 268 462 272
rect 466 268 467 272
rect 481 271 487 272
rect 461 267 467 268
rect 152 264 158 265
rect 142 262 148 263
rect 142 258 143 262
rect 147 258 148 262
rect 142 257 148 258
rect 143 252 145 257
rect 156 255 158 264
rect 465 254 467 267
rect 475 265 477 268
rect 481 267 482 271
rect 486 267 487 271
rect 788 275 794 276
rect 802 275 804 284
rect 812 275 814 284
rect 1114 289 1116 295
rect 1153 289 1155 295
rect 1174 289 1176 295
rect 1207 289 1209 295
rect 1228 289 1230 295
rect 1263 289 1265 295
rect 1284 289 1286 295
rect 1317 289 1319 295
rect 1338 289 1340 295
rect 1383 293 1385 298
rect 788 271 789 275
rect 793 271 794 275
rect 808 274 814 275
rect 788 270 794 271
rect 481 266 487 267
rect 471 264 477 265
rect 471 260 472 264
rect 476 260 477 264
rect 471 259 477 260
rect 472 254 474 259
rect 485 257 487 266
rect 792 257 794 270
rect 802 268 804 271
rect 808 270 809 274
rect 813 270 814 274
rect 1042 272 1044 283
rect 808 269 814 270
rect 798 267 804 268
rect 798 263 799 267
rect 803 263 804 267
rect 798 262 804 263
rect 799 257 801 262
rect 812 260 814 269
rect 1114 271 1116 283
rect 1153 271 1155 283
rect 1174 271 1176 283
rect 1207 271 1209 283
rect 1228 271 1230 283
rect 1263 271 1265 283
rect 1284 271 1286 283
rect 1317 271 1319 283
rect 1338 271 1340 283
rect 1689 305 1695 307
rect 1689 301 1690 305
rect 1694 301 1695 305
rect 1649 299 1653 301
rect 1680 299 1685 301
rect 1689 300 1695 301
rect 1683 293 1685 299
rect 1715 296 1717 317
rect 1728 326 1732 328
rect 1738 327 1762 328
rect 1738 326 1748 327
rect 1747 323 1748 326
rect 1752 326 1762 327
rect 1774 326 1778 328
rect 1752 323 1753 326
rect 1747 322 1753 323
rect 1728 316 1732 318
rect 1738 316 1747 318
rect 1751 317 1760 318
rect 1751 316 1755 317
rect 1754 313 1755 316
rect 1759 315 1760 317
rect 1759 313 1765 315
rect 1783 313 1787 315
rect 1754 312 1760 313
rect 1728 306 1732 308
rect 1738 307 1765 308
rect 1738 306 1747 307
rect 1746 303 1747 306
rect 1751 306 1765 307
rect 1783 306 1787 308
rect 1751 303 1752 306
rect 1746 302 1752 303
rect 1705 294 1717 296
rect 1705 293 1707 294
rect 1683 291 1693 293
rect 1702 291 1707 293
rect 1683 290 1685 291
rect 1668 289 1685 290
rect 1668 285 1669 289
rect 1673 288 1685 289
rect 1673 285 1674 288
rect 1668 284 1674 285
rect 1612 282 1618 283
rect 1612 279 1613 282
rect 1601 278 1613 279
rect 1617 278 1618 282
rect 1601 277 1618 278
rect 1601 276 1603 277
rect 1383 273 1385 276
rect 1395 273 1397 276
rect 1579 274 1584 276
rect 1593 274 1603 276
rect 1579 273 1581 274
rect 156 239 158 243
rect 485 241 487 245
rect 812 244 814 248
rect 1042 250 1044 268
rect 1154 267 1155 271
rect 1175 267 1176 271
rect 1208 267 1209 271
rect 1229 267 1230 271
rect 1264 267 1265 271
rect 1285 267 1286 271
rect 1318 267 1319 271
rect 1339 267 1340 271
rect 1379 272 1385 273
rect 1379 268 1380 272
rect 1384 268 1385 272
rect 1379 267 1385 268
rect 1391 272 1397 273
rect 1391 268 1392 272
rect 1396 268 1397 272
rect 1391 267 1397 268
rect 1042 244 1044 247
rect 1114 249 1116 267
rect 1153 252 1155 267
rect 1174 252 1176 267
rect 1207 252 1209 267
rect 1228 252 1230 267
rect 1263 252 1265 267
rect 1284 252 1286 267
rect 1317 252 1319 267
rect 1338 252 1340 267
rect 1383 264 1385 267
rect 1395 264 1397 267
rect 1569 271 1581 273
rect 1383 249 1385 254
rect 1569 250 1571 271
rect 1601 268 1603 274
rect 1591 266 1597 267
rect 1601 266 1606 268
rect 1633 266 1637 268
rect 1591 262 1592 266
rect 1596 262 1597 266
rect 1591 260 1597 262
rect 1575 258 1579 260
rect 1588 258 1603 260
rect 1601 252 1603 258
rect 1601 250 1606 252
rect 1624 250 1628 252
rect 1114 243 1116 246
rect 1153 243 1155 246
rect 1174 243 1176 246
rect 1207 243 1209 246
rect 1228 243 1230 246
rect 1263 243 1265 246
rect 1284 243 1286 246
rect 1317 243 1319 246
rect 1338 243 1340 246
rect 1395 245 1397 250
rect 1569 248 1579 250
rect 1588 248 1593 250
rect 1597 245 1603 246
rect 1597 242 1598 245
rect 136 230 138 234
rect 143 230 145 234
rect 465 232 467 236
rect 472 232 474 236
rect 792 235 794 239
rect 799 235 801 239
rect 1591 241 1598 242
rect 1602 242 1603 245
rect 1602 241 1606 242
rect 1591 240 1606 241
rect 1624 240 1628 242
rect 1571 238 1576 240
rect 1588 238 1593 240
rect 1118 227 1120 230
rect 1157 227 1159 230
rect 1178 227 1180 230
rect 1211 227 1213 230
rect 1232 227 1234 230
rect 1267 227 1269 230
rect 1288 227 1290 230
rect 1321 227 1323 230
rect 1342 227 1344 230
rect 128 218 130 222
rect 52 210 58 211
rect 42 202 44 207
rect 52 206 53 210
rect 57 206 58 210
rect 52 205 58 206
rect 52 200 54 205
rect 62 200 64 205
rect 113 202 119 203
rect 113 198 114 202
rect 118 198 119 202
rect 113 197 119 198
rect 42 187 44 190
rect 52 187 54 190
rect 42 186 48 187
rect 42 182 43 186
rect 47 182 48 186
rect 52 184 56 187
rect 42 181 48 182
rect 42 173 44 181
rect 54 170 56 184
rect 62 179 64 190
rect 117 188 119 197
rect 164 218 166 222
rect 212 218 214 222
rect 144 209 146 213
rect 154 209 156 213
rect 197 202 203 203
rect 197 198 198 202
rect 202 198 203 202
rect 197 197 203 198
rect 128 188 130 191
rect 144 188 146 191
rect 154 188 156 191
rect 164 188 166 191
rect 117 186 130 188
rect 136 186 146 188
rect 150 187 156 188
rect 61 178 67 179
rect 120 178 122 186
rect 136 182 138 186
rect 150 183 151 187
rect 155 183 156 187
rect 150 182 156 183
rect 160 187 166 188
rect 160 183 161 187
rect 165 183 166 187
rect 201 188 203 197
rect 248 218 250 222
rect 228 209 230 213
rect 238 209 240 213
rect 457 220 459 224
rect 381 212 387 213
rect 284 210 290 211
rect 274 202 276 207
rect 284 206 285 210
rect 289 206 290 210
rect 284 205 290 206
rect 212 188 214 191
rect 228 188 230 191
rect 238 188 240 191
rect 248 188 250 191
rect 284 200 286 205
rect 294 200 296 205
rect 371 204 373 209
rect 381 208 382 212
rect 386 208 387 212
rect 381 207 387 208
rect 381 202 383 207
rect 391 202 393 207
rect 442 204 448 205
rect 442 200 443 204
rect 447 200 448 204
rect 442 199 448 200
rect 201 186 214 188
rect 220 186 230 188
rect 234 187 240 188
rect 160 182 166 183
rect 129 181 138 182
rect 61 174 62 178
rect 66 174 67 178
rect 61 173 67 174
rect 61 170 63 173
rect 42 163 44 167
rect 129 177 130 181
rect 134 177 138 181
rect 154 178 156 182
rect 129 176 138 177
rect 136 173 138 176
rect 146 173 148 178
rect 154 176 158 178
rect 156 173 158 176
rect 163 173 165 182
rect 204 178 206 186
rect 220 182 222 186
rect 234 183 235 187
rect 239 183 240 187
rect 234 182 240 183
rect 244 187 250 188
rect 244 183 245 187
rect 249 183 250 187
rect 244 182 250 183
rect 274 187 276 190
rect 284 187 286 190
rect 274 186 280 187
rect 274 182 275 186
rect 279 182 280 186
rect 284 184 288 187
rect 213 181 222 182
rect 120 166 122 169
rect 120 164 125 166
rect 54 156 56 161
rect 61 156 63 161
rect 123 156 125 164
rect 136 160 138 164
rect 146 156 148 164
rect 213 177 214 181
rect 218 177 222 181
rect 238 178 240 182
rect 213 176 222 177
rect 220 173 222 176
rect 230 173 232 178
rect 238 176 242 178
rect 240 173 242 176
rect 247 173 249 182
rect 274 181 280 182
rect 274 173 276 181
rect 204 166 206 169
rect 204 164 209 166
rect 156 156 158 161
rect 163 156 165 161
rect 123 154 148 156
rect 207 156 209 164
rect 220 160 222 164
rect 230 156 232 164
rect 286 170 288 184
rect 294 179 296 190
rect 371 189 373 192
rect 381 189 383 192
rect 371 188 377 189
rect 371 184 372 188
rect 376 184 377 188
rect 381 186 385 189
rect 371 183 377 184
rect 293 178 299 179
rect 293 174 294 178
rect 298 174 299 178
rect 371 175 373 183
rect 293 173 299 174
rect 293 170 295 173
rect 274 163 276 167
rect 383 172 385 186
rect 391 181 393 192
rect 446 190 448 199
rect 493 220 495 224
rect 541 220 543 224
rect 473 211 475 215
rect 483 211 485 215
rect 526 204 532 205
rect 526 200 527 204
rect 531 200 532 204
rect 526 199 532 200
rect 457 190 459 193
rect 473 190 475 193
rect 483 190 485 193
rect 493 190 495 193
rect 446 188 459 190
rect 465 188 475 190
rect 479 189 485 190
rect 390 180 396 181
rect 449 180 451 188
rect 465 184 467 188
rect 479 185 480 189
rect 484 185 485 189
rect 479 184 485 185
rect 489 189 495 190
rect 489 185 490 189
rect 494 185 495 189
rect 530 190 532 199
rect 577 220 579 224
rect 557 211 559 215
rect 567 211 569 215
rect 784 223 786 227
rect 708 215 714 216
rect 613 212 619 213
rect 603 204 605 209
rect 613 208 614 212
rect 618 208 619 212
rect 613 207 619 208
rect 698 207 700 212
rect 708 211 709 215
rect 713 211 714 215
rect 708 210 714 211
rect 541 190 543 193
rect 557 190 559 193
rect 567 190 569 193
rect 577 190 579 193
rect 613 202 615 207
rect 623 202 625 207
rect 708 205 710 210
rect 718 205 720 210
rect 769 207 775 208
rect 769 203 770 207
rect 774 203 775 207
rect 769 202 775 203
rect 698 192 700 195
rect 708 192 710 195
rect 530 188 543 190
rect 549 188 559 190
rect 563 189 569 190
rect 489 184 495 185
rect 458 183 467 184
rect 390 176 391 180
rect 395 176 396 180
rect 390 175 396 176
rect 390 172 392 175
rect 371 165 373 169
rect 458 179 459 183
rect 463 179 467 183
rect 483 180 485 184
rect 458 178 467 179
rect 465 175 467 178
rect 475 175 477 180
rect 483 178 487 180
rect 485 175 487 178
rect 492 175 494 184
rect 533 180 535 188
rect 549 184 551 188
rect 563 185 564 189
rect 568 185 569 189
rect 563 184 569 185
rect 573 189 579 190
rect 573 185 574 189
rect 578 185 579 189
rect 573 184 579 185
rect 603 189 605 192
rect 613 189 615 192
rect 603 188 609 189
rect 603 184 604 188
rect 608 184 609 188
rect 613 186 617 189
rect 542 183 551 184
rect 449 168 451 171
rect 449 166 454 168
rect 240 156 242 161
rect 247 156 249 161
rect 207 154 232 156
rect 286 156 288 161
rect 293 156 295 161
rect 383 158 385 163
rect 390 158 392 163
rect 452 158 454 166
rect 465 162 467 166
rect 475 158 477 166
rect 542 179 543 183
rect 547 179 551 183
rect 567 180 569 184
rect 542 178 551 179
rect 549 175 551 178
rect 559 175 561 180
rect 567 178 571 180
rect 569 175 571 178
rect 576 175 578 184
rect 603 183 609 184
rect 603 175 605 183
rect 533 168 535 171
rect 533 166 538 168
rect 485 158 487 163
rect 492 158 494 163
rect 452 156 477 158
rect 536 158 538 166
rect 549 162 551 166
rect 559 158 561 166
rect 615 172 617 186
rect 623 181 625 192
rect 698 191 704 192
rect 698 187 699 191
rect 703 187 704 191
rect 708 189 712 192
rect 698 186 704 187
rect 622 180 628 181
rect 622 176 623 180
rect 627 176 628 180
rect 698 178 700 186
rect 622 175 628 176
rect 622 172 624 175
rect 710 175 712 189
rect 718 184 720 195
rect 773 193 775 202
rect 820 223 822 227
rect 868 223 870 227
rect 800 214 802 218
rect 810 214 812 218
rect 853 207 859 208
rect 853 203 854 207
rect 858 203 859 207
rect 853 202 859 203
rect 784 193 786 196
rect 800 193 802 196
rect 810 193 812 196
rect 820 193 822 196
rect 773 191 786 193
rect 792 191 802 193
rect 806 192 812 193
rect 717 183 723 184
rect 776 183 778 191
rect 792 187 794 191
rect 806 188 807 192
rect 811 188 812 192
rect 806 187 812 188
rect 816 192 822 193
rect 816 188 817 192
rect 821 188 822 192
rect 857 193 859 202
rect 904 223 906 227
rect 884 214 886 218
rect 894 214 896 218
rect 940 215 946 216
rect 930 207 932 212
rect 940 211 941 215
rect 945 211 946 215
rect 940 210 946 211
rect 868 193 870 196
rect 884 193 886 196
rect 894 193 896 196
rect 904 193 906 196
rect 940 205 942 210
rect 950 205 952 210
rect 1118 206 1120 224
rect 1384 225 1386 230
rect 1396 229 1398 234
rect 1597 235 1603 236
rect 1597 233 1598 235
rect 1571 231 1576 233
rect 1588 231 1598 233
rect 1602 232 1603 235
rect 1602 231 1606 232
rect 1597 230 1606 231
rect 1633 230 1637 232
rect 1157 206 1159 221
rect 1178 206 1180 221
rect 1211 206 1213 221
rect 1232 206 1234 221
rect 1267 206 1269 221
rect 1288 206 1290 221
rect 1321 206 1323 221
rect 1342 206 1344 221
rect 1692 237 1698 238
rect 1692 235 1693 237
rect 1666 233 1671 235
rect 1681 233 1693 235
rect 1697 234 1698 237
rect 1697 233 1701 234
rect 1692 232 1701 233
rect 1710 232 1715 234
rect 1660 228 1666 229
rect 1660 224 1661 228
rect 1665 225 1666 228
rect 1684 225 1701 227
rect 1710 225 1715 227
rect 1665 224 1671 225
rect 1660 223 1671 224
rect 1681 223 1687 225
rect 1384 212 1386 215
rect 1396 212 1398 215
rect 1380 211 1386 212
rect 1380 207 1381 211
rect 1385 207 1386 211
rect 1380 206 1386 207
rect 1392 211 1398 212
rect 1392 207 1393 211
rect 1397 207 1398 211
rect 1392 206 1398 207
rect 1684 218 1690 219
rect 1684 215 1685 218
rect 1664 213 1669 215
rect 1681 214 1685 215
rect 1689 215 1690 218
rect 1689 214 1698 215
rect 1681 213 1698 214
rect 1704 213 1708 215
rect 1158 202 1159 206
rect 1179 202 1180 206
rect 1212 202 1213 206
rect 1233 202 1234 206
rect 1268 202 1269 206
rect 1289 202 1290 206
rect 1322 202 1323 206
rect 1343 202 1344 206
rect 1384 203 1386 206
rect 1396 203 1398 206
rect 1578 204 1582 206
rect 1588 205 1605 206
rect 1588 204 1597 205
rect 857 191 870 193
rect 876 191 886 193
rect 890 192 896 193
rect 816 187 822 188
rect 785 186 794 187
rect 717 179 718 183
rect 722 179 723 183
rect 717 178 723 179
rect 717 175 719 178
rect 603 165 605 169
rect 698 168 700 172
rect 785 182 786 186
rect 790 182 794 186
rect 810 183 812 187
rect 785 181 794 182
rect 792 178 794 181
rect 802 178 804 183
rect 810 181 814 183
rect 812 178 814 181
rect 819 178 821 187
rect 860 183 862 191
rect 876 187 878 191
rect 890 188 891 192
rect 895 188 896 192
rect 890 187 896 188
rect 900 192 906 193
rect 900 188 901 192
rect 905 188 906 192
rect 900 187 906 188
rect 930 192 932 195
rect 940 192 942 195
rect 930 191 936 192
rect 930 187 931 191
rect 935 187 936 191
rect 940 189 944 192
rect 869 186 878 187
rect 776 171 778 174
rect 776 169 781 171
rect 569 158 571 163
rect 576 158 578 163
rect 536 156 561 158
rect 615 158 617 163
rect 622 158 624 163
rect 710 161 712 166
rect 717 161 719 166
rect 779 161 781 169
rect 792 165 794 169
rect 802 161 804 169
rect 869 182 870 186
rect 874 182 878 186
rect 894 183 896 187
rect 869 181 878 182
rect 876 178 878 181
rect 886 178 888 183
rect 894 181 898 183
rect 896 178 898 181
rect 903 178 905 187
rect 930 186 936 187
rect 930 178 932 186
rect 860 171 862 174
rect 860 169 865 171
rect 812 161 814 166
rect 819 161 821 166
rect 779 159 804 161
rect 863 161 865 169
rect 876 165 878 169
rect 886 161 888 169
rect 942 175 944 189
rect 950 184 952 195
rect 1118 190 1120 202
rect 1157 190 1159 202
rect 1178 190 1180 202
rect 1211 190 1213 202
rect 1232 190 1234 202
rect 1267 190 1269 202
rect 1288 190 1290 202
rect 1321 190 1323 202
rect 1342 190 1344 202
rect 949 183 955 184
rect 949 179 950 183
rect 954 179 955 183
rect 949 178 955 179
rect 1118 178 1120 184
rect 1157 178 1159 184
rect 1178 178 1180 184
rect 1211 178 1213 184
rect 1232 178 1234 184
rect 1267 178 1269 184
rect 1288 178 1290 184
rect 1321 178 1323 184
rect 1342 178 1344 184
rect 1384 181 1386 186
rect 949 175 951 178
rect 930 168 932 172
rect 1596 201 1597 204
rect 1601 204 1605 205
rect 1617 204 1622 206
rect 1601 201 1602 204
rect 1596 200 1602 201
rect 1599 194 1605 196
rect 1615 195 1626 196
rect 1615 194 1621 195
rect 1571 192 1576 194
rect 1585 192 1602 194
rect 1620 191 1621 194
rect 1625 191 1626 195
rect 1620 190 1626 191
rect 1571 185 1576 187
rect 1585 186 1594 187
rect 1585 185 1589 186
rect 1588 182 1589 185
rect 1593 184 1605 186
rect 1615 184 1620 186
rect 1593 182 1594 184
rect 1588 181 1594 182
rect 1396 171 1398 175
rect 896 161 898 166
rect 903 161 905 166
rect 863 159 888 161
rect 942 161 944 166
rect 949 161 951 166
rect 1395 164 1397 168
rect 1383 153 1385 158
rect 135 139 137 143
rect 145 139 147 143
rect 155 139 157 143
rect 464 141 466 145
rect 474 141 476 145
rect 484 141 486 145
rect 791 144 793 148
rect 801 144 803 148
rect 811 144 813 148
rect 1041 147 1043 149
rect 1113 147 1115 153
rect 1152 147 1154 153
rect 1173 147 1175 153
rect 1206 147 1208 153
rect 1227 147 1229 153
rect 1262 147 1264 153
rect 1283 147 1285 153
rect 1316 147 1318 153
rect 1337 147 1339 153
rect 135 125 137 133
rect 131 124 137 125
rect 145 124 147 133
rect 155 124 157 133
rect 464 127 466 135
rect 131 120 132 124
rect 136 120 137 124
rect 151 123 157 124
rect 131 119 137 120
rect 135 106 137 119
rect 145 117 147 120
rect 151 119 152 123
rect 156 119 157 123
rect 460 126 466 127
rect 474 126 476 135
rect 484 126 486 135
rect 791 130 793 138
rect 460 122 461 126
rect 465 122 466 126
rect 480 125 486 126
rect 460 121 466 122
rect 151 118 157 119
rect 141 116 147 117
rect 141 112 142 116
rect 146 112 147 116
rect 141 111 147 112
rect 142 106 144 111
rect 155 109 157 118
rect 464 108 466 121
rect 474 119 476 122
rect 480 121 481 125
rect 485 121 486 125
rect 787 129 793 130
rect 801 129 803 138
rect 811 129 813 138
rect 1041 130 1043 141
rect 787 125 788 129
rect 792 125 793 129
rect 807 128 813 129
rect 787 124 793 125
rect 480 120 486 121
rect 470 118 476 119
rect 470 114 471 118
rect 475 114 476 118
rect 470 113 476 114
rect 471 108 473 113
rect 484 111 486 120
rect 791 111 793 124
rect 801 122 803 125
rect 807 124 808 128
rect 812 124 813 128
rect 1113 129 1115 141
rect 1152 129 1154 141
rect 1173 129 1175 141
rect 1206 129 1208 141
rect 1227 129 1229 141
rect 1262 129 1264 141
rect 1283 129 1285 141
rect 1316 129 1318 141
rect 1337 129 1339 141
rect 1383 133 1385 136
rect 1395 133 1397 136
rect 807 123 813 124
rect 797 121 803 122
rect 797 117 798 121
rect 802 117 803 121
rect 797 116 803 117
rect 798 111 800 116
rect 811 114 813 123
rect 155 93 157 97
rect 484 95 486 99
rect 1041 108 1043 126
rect 1153 125 1154 129
rect 1174 125 1175 129
rect 1207 125 1208 129
rect 1228 125 1229 129
rect 1263 125 1264 129
rect 1284 125 1285 129
rect 1317 125 1318 129
rect 1338 125 1339 129
rect 1379 132 1385 133
rect 1379 128 1380 132
rect 1384 128 1385 132
rect 1379 127 1385 128
rect 1391 132 1397 133
rect 1391 128 1392 132
rect 1396 128 1397 132
rect 1391 127 1397 128
rect 1041 102 1043 105
rect 1113 107 1115 125
rect 1152 110 1154 125
rect 1173 110 1175 125
rect 1206 110 1208 125
rect 1227 110 1229 125
rect 1262 110 1264 125
rect 1283 110 1285 125
rect 1316 110 1318 125
rect 1337 110 1339 125
rect 1383 124 1385 127
rect 1395 124 1397 127
rect 1383 109 1385 114
rect 811 98 813 102
rect 1113 101 1115 104
rect 1152 101 1154 104
rect 1173 101 1175 104
rect 1206 101 1208 104
rect 1227 101 1229 104
rect 1262 101 1264 104
rect 1283 101 1285 104
rect 1316 101 1318 104
rect 1337 101 1339 104
rect 1395 105 1397 110
rect 1694 109 1700 110
rect 1694 107 1695 109
rect 1668 105 1673 107
rect 1683 105 1695 107
rect 1699 106 1700 109
rect 1699 105 1703 106
rect 1694 104 1703 105
rect 1712 104 1717 106
rect 135 84 137 88
rect 142 84 144 88
rect 464 86 466 90
rect 471 86 473 90
rect 791 89 793 93
rect 798 89 800 93
rect 1662 100 1668 101
rect 1662 96 1663 100
rect 1667 97 1668 100
rect 1686 97 1703 99
rect 1712 97 1717 99
rect 1667 96 1673 97
rect 1662 95 1673 96
rect 1683 95 1689 97
rect 1117 85 1119 88
rect 1156 85 1158 88
rect 1177 85 1179 88
rect 1210 85 1212 88
rect 1231 85 1233 88
rect 1266 85 1268 88
rect 1287 85 1289 88
rect 1320 85 1322 88
rect 1341 85 1343 88
rect 336 61 338 65
rect 346 63 348 68
rect 356 63 358 68
rect 429 61 431 65
rect 439 63 441 68
rect 449 63 451 68
rect 336 39 338 43
rect 346 39 348 50
rect 356 47 358 50
rect 356 46 362 47
rect 356 42 357 46
rect 361 42 362 46
rect 516 61 518 65
rect 526 63 528 68
rect 536 63 538 68
rect 1117 64 1119 82
rect 1156 64 1158 79
rect 1177 64 1179 79
rect 1210 64 1212 79
rect 1231 64 1233 79
rect 1266 64 1268 79
rect 1287 64 1289 79
rect 1320 64 1322 79
rect 1341 64 1343 79
rect 1686 90 1692 91
rect 1686 87 1687 90
rect 1666 85 1671 87
rect 1683 86 1687 87
rect 1691 87 1692 90
rect 1691 86 1700 87
rect 1683 85 1700 86
rect 1706 85 1710 87
rect 1580 76 1584 78
rect 1590 77 1607 78
rect 1590 76 1599 77
rect 1598 73 1599 76
rect 1603 76 1607 77
rect 1619 76 1624 78
rect 1603 73 1604 76
rect 1598 72 1604 73
rect 1601 66 1607 68
rect 1617 67 1628 68
rect 1617 66 1623 67
rect 1573 64 1578 66
rect 1587 64 1604 66
rect 356 41 362 42
rect 336 38 342 39
rect 336 34 337 38
rect 341 34 342 38
rect 336 33 342 34
rect 346 38 352 39
rect 346 34 347 38
rect 351 34 352 38
rect 346 33 352 34
rect 336 28 338 33
rect 349 28 351 33
rect 356 28 358 41
rect 429 39 431 43
rect 439 39 441 50
rect 449 47 451 50
rect 449 46 455 47
rect 449 42 450 46
rect 454 42 455 46
rect 1157 60 1158 64
rect 1178 60 1179 64
rect 1211 60 1212 64
rect 1232 60 1233 64
rect 1267 60 1268 64
rect 1288 60 1289 64
rect 1321 60 1322 64
rect 1342 60 1343 64
rect 449 41 455 42
rect 429 38 435 39
rect 429 34 430 38
rect 434 34 435 38
rect 429 33 435 34
rect 439 38 445 39
rect 439 34 440 38
rect 444 34 445 38
rect 439 33 445 34
rect 429 28 431 33
rect 442 28 444 33
rect 449 28 451 41
rect 516 39 518 43
rect 526 39 528 50
rect 536 47 538 50
rect 1117 48 1119 60
rect 1156 48 1158 60
rect 1177 48 1179 60
rect 1210 48 1212 60
rect 1231 48 1233 60
rect 1266 48 1268 60
rect 1287 48 1289 60
rect 1320 48 1322 60
rect 1341 48 1343 60
rect 1622 63 1623 66
rect 1627 63 1628 67
rect 1622 62 1628 63
rect 1573 57 1578 59
rect 1587 58 1596 59
rect 1587 57 1591 58
rect 1590 54 1591 57
rect 1595 56 1607 58
rect 1617 56 1622 58
rect 1595 54 1596 56
rect 1590 53 1596 54
rect 1651 59 1655 61
rect 1682 60 1691 61
rect 1682 59 1686 60
rect 1685 56 1686 59
rect 1690 58 1700 60
rect 1712 58 1717 60
rect 1690 56 1691 58
rect 1685 55 1691 56
rect 1695 51 1700 53
rect 1712 51 1717 53
rect 1660 49 1664 51
rect 1682 50 1697 51
rect 1682 49 1686 50
rect 536 46 542 47
rect 536 42 537 46
rect 541 42 542 46
rect 1685 46 1686 49
rect 1690 49 1697 50
rect 1690 46 1691 49
rect 1685 45 1691 46
rect 536 41 542 42
rect 516 38 522 39
rect 516 34 517 38
rect 521 34 522 38
rect 516 33 522 34
rect 526 38 532 39
rect 526 34 527 38
rect 531 34 532 38
rect 526 33 532 34
rect 516 28 518 33
rect 529 28 531 33
rect 536 28 538 41
rect 1117 36 1119 42
rect 1156 36 1158 42
rect 1177 36 1179 42
rect 1210 36 1212 42
rect 1231 36 1233 42
rect 1266 36 1268 42
rect 1287 36 1289 42
rect 1320 36 1322 42
rect 1341 36 1343 42
rect 1695 41 1700 43
rect 1709 41 1719 43
rect 1660 39 1664 41
rect 1682 39 1687 41
rect 1685 33 1687 39
rect 1685 31 1700 33
rect 1709 31 1713 33
rect 336 15 338 19
rect 349 12 351 17
rect 356 12 358 17
rect 429 15 431 19
rect 442 12 444 17
rect 449 12 451 17
rect 516 15 518 19
rect 1691 29 1697 31
rect 1691 25 1692 29
rect 1696 25 1697 29
rect 1651 23 1655 25
rect 1682 23 1687 25
rect 1691 24 1697 25
rect 529 12 531 17
rect 536 12 538 17
rect 1685 17 1687 23
rect 1717 20 1719 41
rect 1707 18 1719 20
rect 1707 17 1709 18
rect 1685 15 1695 17
rect 1704 15 1709 17
rect 1685 14 1687 15
rect 1670 13 1687 14
rect 1670 9 1671 13
rect 1675 12 1687 13
rect 1675 9 1676 12
rect 1670 8 1676 9
rect 1614 6 1620 7
rect 1614 3 1615 6
rect 1603 2 1615 3
rect 1619 2 1620 6
rect 1603 1 1620 2
rect 1603 0 1605 1
rect 1581 -2 1586 0
rect 1595 -2 1605 0
rect 1581 -3 1583 -2
rect 1571 -5 1583 -3
rect 1536 -12 1542 -11
rect 1536 -15 1537 -12
rect 1501 -17 1505 -15
rect 1523 -16 1537 -15
rect 1541 -15 1542 -12
rect 1541 -16 1550 -15
rect 1523 -17 1550 -16
rect 1556 -17 1560 -15
rect 1528 -22 1534 -21
rect 1501 -24 1505 -22
rect 1523 -24 1529 -22
rect 1528 -26 1529 -24
rect 1533 -25 1534 -22
rect 1533 -26 1537 -25
rect 1528 -27 1537 -26
rect 1541 -27 1550 -25
rect 1556 -27 1560 -25
rect 1535 -32 1541 -31
rect 1535 -35 1536 -32
rect 1510 -37 1514 -35
rect 1526 -36 1536 -35
rect 1540 -35 1541 -32
rect 1540 -36 1550 -35
rect 1526 -37 1550 -36
rect 1556 -37 1560 -35
rect 1571 -26 1573 -5
rect 1603 -8 1605 -2
rect 1593 -10 1599 -9
rect 1603 -10 1608 -8
rect 1635 -10 1639 -8
rect 1593 -14 1594 -10
rect 1598 -14 1599 -10
rect 1593 -16 1599 -14
rect 1577 -18 1581 -16
rect 1590 -18 1605 -16
rect 1603 -24 1605 -18
rect 1603 -26 1608 -24
rect 1626 -26 1630 -24
rect 1651 -25 1655 -23
rect 1682 -24 1691 -23
rect 1682 -25 1686 -24
rect 1571 -28 1581 -26
rect 1590 -28 1595 -26
rect 1599 -31 1605 -30
rect 1599 -34 1600 -31
rect 1593 -35 1600 -34
rect 1604 -34 1605 -31
rect 1685 -28 1686 -25
rect 1690 -26 1700 -24
rect 1712 -26 1717 -24
rect 1690 -28 1691 -26
rect 1685 -29 1691 -28
rect 1695 -33 1700 -31
rect 1712 -33 1717 -31
rect 1604 -35 1608 -34
rect 1593 -36 1608 -35
rect 1626 -36 1630 -34
rect 1660 -35 1664 -33
rect 1682 -34 1697 -33
rect 1682 -35 1686 -34
rect 1573 -38 1578 -36
rect 1590 -38 1595 -36
rect 1599 -41 1605 -40
rect 1599 -43 1600 -41
rect 1573 -45 1578 -43
rect 1590 -45 1600 -43
rect 1604 -44 1605 -41
rect 1685 -38 1686 -35
rect 1690 -35 1697 -34
rect 1690 -38 1691 -35
rect 1685 -39 1691 -38
rect 1695 -43 1700 -41
rect 1709 -43 1719 -41
rect 1604 -45 1608 -44
rect 1599 -46 1608 -45
rect 1635 -46 1639 -44
rect 1660 -45 1664 -43
rect 1682 -45 1687 -43
rect 1685 -51 1687 -45
rect 1685 -53 1700 -51
rect 1709 -53 1713 -51
rect 132 -70 134 -65
rect 139 -70 141 -65
rect 152 -72 154 -68
rect 219 -70 221 -65
rect 226 -70 228 -65
rect 239 -72 241 -68
rect 312 -70 314 -65
rect 319 -70 321 -65
rect 332 -72 334 -68
rect 552 -70 554 -66
rect 565 -68 567 -63
rect 572 -68 574 -63
rect 645 -70 647 -66
rect 658 -68 660 -63
rect 665 -68 667 -63
rect 1691 -55 1697 -53
rect 1691 -59 1692 -55
rect 1696 -59 1697 -55
rect 1651 -61 1655 -59
rect 1682 -61 1687 -59
rect 1691 -60 1697 -59
rect 732 -70 734 -66
rect 745 -68 747 -63
rect 752 -68 754 -63
rect 1685 -67 1687 -61
rect 1717 -64 1719 -43
rect 1730 -34 1734 -32
rect 1740 -33 1764 -32
rect 1740 -34 1750 -33
rect 1749 -37 1750 -34
rect 1754 -34 1764 -33
rect 1776 -34 1780 -32
rect 1754 -37 1755 -34
rect 1749 -38 1755 -37
rect 1730 -44 1734 -42
rect 1740 -44 1749 -42
rect 1753 -43 1762 -42
rect 1753 -44 1757 -43
rect 1756 -47 1757 -44
rect 1761 -45 1762 -43
rect 1761 -47 1767 -45
rect 1785 -47 1789 -45
rect 1756 -48 1762 -47
rect 1730 -54 1734 -52
rect 1740 -53 1767 -52
rect 1740 -54 1749 -53
rect 1748 -57 1749 -54
rect 1753 -54 1767 -53
rect 1785 -54 1789 -52
rect 1753 -57 1754 -54
rect 1748 -58 1754 -57
rect 1707 -66 1719 -64
rect 1707 -67 1709 -66
rect 1685 -69 1695 -67
rect 1704 -69 1709 -67
rect 1685 -70 1687 -69
rect 1670 -71 1687 -70
rect 1063 -77 1065 -75
rect 132 -94 134 -81
rect 139 -86 141 -81
rect 152 -86 154 -81
rect 138 -87 144 -86
rect 138 -91 139 -87
rect 143 -91 144 -87
rect 138 -92 144 -91
rect 148 -87 154 -86
rect 148 -91 149 -87
rect 153 -91 154 -87
rect 148 -92 154 -91
rect 128 -95 134 -94
rect 128 -99 129 -95
rect 133 -99 134 -95
rect 128 -100 134 -99
rect 132 -103 134 -100
rect 142 -103 144 -92
rect 152 -96 154 -92
rect 219 -94 221 -81
rect 226 -86 228 -81
rect 239 -86 241 -81
rect 225 -87 231 -86
rect 225 -91 226 -87
rect 230 -91 231 -87
rect 225 -92 231 -91
rect 235 -87 241 -86
rect 235 -91 236 -87
rect 240 -91 241 -87
rect 235 -92 241 -91
rect 215 -95 221 -94
rect 215 -99 216 -95
rect 220 -99 221 -95
rect 215 -100 221 -99
rect 219 -103 221 -100
rect 229 -103 231 -92
rect 239 -96 241 -92
rect 312 -94 314 -81
rect 319 -86 321 -81
rect 332 -86 334 -81
rect 318 -87 324 -86
rect 318 -91 319 -87
rect 323 -91 324 -87
rect 318 -92 324 -91
rect 328 -87 334 -86
rect 328 -91 329 -87
rect 333 -91 334 -87
rect 328 -92 334 -91
rect 308 -95 314 -94
rect 132 -121 134 -116
rect 142 -121 144 -116
rect 152 -118 154 -114
rect 308 -99 309 -95
rect 313 -99 314 -95
rect 308 -100 314 -99
rect 312 -103 314 -100
rect 322 -103 324 -92
rect 332 -96 334 -92
rect 552 -84 554 -79
rect 565 -84 567 -79
rect 552 -85 558 -84
rect 552 -89 553 -85
rect 557 -89 558 -85
rect 552 -90 558 -89
rect 562 -85 568 -84
rect 562 -89 563 -85
rect 567 -89 568 -85
rect 562 -90 568 -89
rect 552 -94 554 -90
rect 219 -121 221 -116
rect 229 -121 231 -116
rect 239 -118 241 -114
rect 562 -101 564 -90
rect 572 -92 574 -79
rect 645 -84 647 -79
rect 658 -84 660 -79
rect 645 -85 651 -84
rect 645 -89 646 -85
rect 650 -89 651 -85
rect 645 -90 651 -89
rect 655 -85 661 -84
rect 655 -89 656 -85
rect 660 -89 661 -85
rect 655 -90 661 -89
rect 572 -93 578 -92
rect 572 -97 573 -93
rect 577 -97 578 -93
rect 645 -94 647 -90
rect 572 -98 578 -97
rect 572 -101 574 -98
rect 312 -121 314 -116
rect 322 -121 324 -116
rect 332 -118 334 -114
rect 552 -116 554 -112
rect 655 -101 657 -90
rect 665 -92 667 -79
rect 732 -84 734 -79
rect 745 -84 747 -79
rect 732 -85 738 -84
rect 732 -89 733 -85
rect 737 -89 738 -85
rect 732 -90 738 -89
rect 742 -85 748 -84
rect 742 -89 743 -85
rect 747 -89 748 -85
rect 742 -90 748 -89
rect 665 -93 671 -92
rect 665 -97 666 -93
rect 670 -97 671 -93
rect 732 -94 734 -90
rect 665 -98 671 -97
rect 665 -101 667 -98
rect 562 -119 564 -114
rect 572 -119 574 -114
rect 645 -116 647 -112
rect 742 -101 744 -90
rect 752 -92 754 -79
rect 1135 -77 1137 -71
rect 1174 -77 1176 -71
rect 1195 -77 1197 -71
rect 1228 -77 1230 -71
rect 1249 -77 1251 -71
rect 1284 -77 1286 -71
rect 1305 -77 1307 -71
rect 1338 -77 1340 -71
rect 1359 -77 1361 -71
rect 1670 -75 1671 -71
rect 1675 -72 1687 -71
rect 1675 -75 1676 -72
rect 1670 -76 1676 -75
rect 752 -93 758 -92
rect 752 -97 753 -93
rect 757 -97 758 -93
rect 1063 -94 1065 -83
rect 752 -98 758 -97
rect 1135 -95 1137 -83
rect 1174 -95 1176 -83
rect 1195 -95 1197 -83
rect 1228 -95 1230 -83
rect 1249 -95 1251 -83
rect 1284 -95 1286 -83
rect 1305 -95 1307 -83
rect 1338 -95 1340 -83
rect 1359 -95 1361 -83
rect 1614 -78 1620 -77
rect 1614 -81 1615 -78
rect 1603 -82 1615 -81
rect 1619 -82 1620 -78
rect 1603 -83 1620 -82
rect 1603 -84 1605 -83
rect 1581 -86 1586 -84
rect 1595 -86 1605 -84
rect 1581 -87 1583 -86
rect 752 -101 754 -98
rect 655 -119 657 -114
rect 665 -119 667 -114
rect 732 -116 734 -112
rect 742 -119 744 -114
rect 752 -119 754 -114
rect 1063 -116 1065 -98
rect 1175 -99 1176 -95
rect 1196 -99 1197 -95
rect 1229 -99 1230 -95
rect 1250 -99 1251 -95
rect 1285 -99 1286 -95
rect 1306 -99 1307 -95
rect 1339 -99 1340 -95
rect 1360 -99 1361 -95
rect 1063 -122 1065 -119
rect 1135 -117 1137 -99
rect 1174 -114 1176 -99
rect 1195 -114 1197 -99
rect 1228 -114 1230 -99
rect 1249 -114 1251 -99
rect 1284 -114 1286 -99
rect 1305 -114 1307 -99
rect 1338 -114 1340 -99
rect 1359 -114 1361 -99
rect 1571 -89 1583 -87
rect 1571 -110 1573 -89
rect 1603 -92 1605 -86
rect 1593 -94 1599 -93
rect 1603 -94 1608 -92
rect 1635 -94 1639 -92
rect 1593 -98 1594 -94
rect 1598 -98 1599 -94
rect 1593 -100 1599 -98
rect 1577 -102 1581 -100
rect 1590 -102 1605 -100
rect 1603 -108 1605 -102
rect 1603 -110 1608 -108
rect 1626 -110 1630 -108
rect 1571 -112 1581 -110
rect 1590 -112 1595 -110
rect 1599 -115 1605 -114
rect 1599 -118 1600 -115
rect 1593 -119 1600 -118
rect 1604 -118 1605 -115
rect 1604 -119 1608 -118
rect 1593 -120 1608 -119
rect 1626 -120 1630 -118
rect 1135 -123 1137 -120
rect 1174 -123 1176 -120
rect 1195 -123 1197 -120
rect 1228 -123 1230 -120
rect 1249 -123 1251 -120
rect 1284 -123 1286 -120
rect 1305 -123 1307 -120
rect 1338 -123 1340 -120
rect 1359 -123 1361 -120
rect 1573 -122 1578 -120
rect 1590 -122 1595 -120
rect 1599 -125 1605 -124
rect 1599 -127 1600 -125
rect 1573 -129 1578 -127
rect 1590 -129 1600 -127
rect 1604 -128 1605 -125
rect 1604 -129 1608 -128
rect 1599 -130 1608 -129
rect 1635 -130 1639 -128
rect 140 -142 142 -138
rect 64 -150 70 -149
rect 54 -158 56 -153
rect 64 -154 65 -150
rect 69 -154 70 -150
rect 64 -155 70 -154
rect 64 -160 66 -155
rect 74 -160 76 -155
rect 125 -158 131 -157
rect 125 -162 126 -158
rect 130 -162 131 -158
rect 125 -163 131 -162
rect 54 -173 56 -170
rect 64 -173 66 -170
rect 54 -174 60 -173
rect 54 -178 55 -174
rect 59 -178 60 -174
rect 64 -176 68 -173
rect 54 -179 60 -178
rect 54 -187 56 -179
rect 66 -190 68 -176
rect 74 -181 76 -170
rect 129 -172 131 -163
rect 176 -142 178 -138
rect 224 -142 226 -138
rect 156 -151 158 -147
rect 166 -151 168 -147
rect 209 -158 215 -157
rect 209 -162 210 -158
rect 214 -162 215 -158
rect 209 -163 215 -162
rect 140 -172 142 -169
rect 156 -172 158 -169
rect 166 -172 168 -169
rect 176 -172 178 -169
rect 129 -174 142 -172
rect 148 -174 158 -172
rect 162 -173 168 -172
rect 73 -182 79 -181
rect 132 -182 134 -174
rect 148 -178 150 -174
rect 162 -177 163 -173
rect 167 -177 168 -173
rect 162 -178 168 -177
rect 172 -173 178 -172
rect 172 -177 173 -173
rect 177 -177 178 -173
rect 213 -172 215 -163
rect 260 -142 262 -138
rect 240 -151 242 -147
rect 250 -151 252 -147
rect 469 -140 471 -136
rect 393 -148 399 -147
rect 296 -150 302 -149
rect 286 -158 288 -153
rect 296 -154 297 -150
rect 301 -154 302 -150
rect 296 -155 302 -154
rect 224 -172 226 -169
rect 240 -172 242 -169
rect 250 -172 252 -169
rect 260 -172 262 -169
rect 296 -160 298 -155
rect 306 -160 308 -155
rect 383 -156 385 -151
rect 393 -152 394 -148
rect 398 -152 399 -148
rect 393 -153 399 -152
rect 393 -158 395 -153
rect 403 -158 405 -153
rect 454 -156 460 -155
rect 454 -160 455 -156
rect 459 -160 460 -156
rect 454 -161 460 -160
rect 213 -174 226 -172
rect 232 -174 242 -172
rect 246 -173 252 -172
rect 172 -178 178 -177
rect 141 -179 150 -178
rect 73 -186 74 -182
rect 78 -186 79 -182
rect 73 -187 79 -186
rect 73 -190 75 -187
rect 54 -197 56 -193
rect 141 -183 142 -179
rect 146 -183 150 -179
rect 166 -182 168 -178
rect 141 -184 150 -183
rect 148 -187 150 -184
rect 158 -187 160 -182
rect 166 -184 170 -182
rect 168 -187 170 -184
rect 175 -187 177 -178
rect 216 -182 218 -174
rect 232 -178 234 -174
rect 246 -177 247 -173
rect 251 -177 252 -173
rect 246 -178 252 -177
rect 256 -173 262 -172
rect 256 -177 257 -173
rect 261 -177 262 -173
rect 256 -178 262 -177
rect 286 -173 288 -170
rect 296 -173 298 -170
rect 286 -174 292 -173
rect 286 -178 287 -174
rect 291 -178 292 -174
rect 296 -176 300 -173
rect 225 -179 234 -178
rect 132 -194 134 -191
rect 132 -196 137 -194
rect 66 -204 68 -199
rect 73 -204 75 -199
rect 135 -204 137 -196
rect 148 -200 150 -196
rect 158 -204 160 -196
rect 225 -183 226 -179
rect 230 -183 234 -179
rect 250 -182 252 -178
rect 225 -184 234 -183
rect 232 -187 234 -184
rect 242 -187 244 -182
rect 250 -184 254 -182
rect 252 -187 254 -184
rect 259 -187 261 -178
rect 286 -179 292 -178
rect 286 -187 288 -179
rect 216 -194 218 -191
rect 216 -196 221 -194
rect 168 -204 170 -199
rect 175 -204 177 -199
rect 135 -206 160 -204
rect 219 -204 221 -196
rect 232 -200 234 -196
rect 242 -204 244 -196
rect 298 -190 300 -176
rect 306 -181 308 -170
rect 383 -171 385 -168
rect 393 -171 395 -168
rect 383 -172 389 -171
rect 383 -176 384 -172
rect 388 -176 389 -172
rect 393 -174 397 -171
rect 383 -177 389 -176
rect 305 -182 311 -181
rect 305 -186 306 -182
rect 310 -186 311 -182
rect 383 -185 385 -177
rect 305 -187 311 -186
rect 305 -190 307 -187
rect 286 -197 288 -193
rect 395 -188 397 -174
rect 403 -179 405 -168
rect 458 -170 460 -161
rect 505 -140 507 -136
rect 553 -140 555 -136
rect 485 -149 487 -145
rect 495 -149 497 -145
rect 538 -156 544 -155
rect 538 -160 539 -156
rect 543 -160 544 -156
rect 538 -161 544 -160
rect 469 -170 471 -167
rect 485 -170 487 -167
rect 495 -170 497 -167
rect 505 -170 507 -167
rect 458 -172 471 -170
rect 477 -172 487 -170
rect 491 -171 497 -170
rect 402 -180 408 -179
rect 461 -180 463 -172
rect 477 -176 479 -172
rect 491 -175 492 -171
rect 496 -175 497 -171
rect 491 -176 497 -175
rect 501 -171 507 -170
rect 501 -175 502 -171
rect 506 -175 507 -171
rect 542 -170 544 -161
rect 589 -140 591 -136
rect 569 -149 571 -145
rect 579 -149 581 -145
rect 796 -137 798 -133
rect 720 -145 726 -144
rect 625 -148 631 -147
rect 615 -156 617 -151
rect 625 -152 626 -148
rect 630 -152 631 -148
rect 625 -153 631 -152
rect 710 -153 712 -148
rect 720 -149 721 -145
rect 725 -149 726 -145
rect 720 -150 726 -149
rect 553 -170 555 -167
rect 569 -170 571 -167
rect 579 -170 581 -167
rect 589 -170 591 -167
rect 625 -158 627 -153
rect 635 -158 637 -153
rect 720 -155 722 -150
rect 730 -155 732 -150
rect 781 -153 787 -152
rect 781 -157 782 -153
rect 786 -157 787 -153
rect 781 -158 787 -157
rect 710 -168 712 -165
rect 720 -168 722 -165
rect 542 -172 555 -170
rect 561 -172 571 -170
rect 575 -171 581 -170
rect 501 -176 507 -175
rect 470 -177 479 -176
rect 402 -184 403 -180
rect 407 -184 408 -180
rect 402 -185 408 -184
rect 402 -188 404 -185
rect 383 -195 385 -191
rect 470 -181 471 -177
rect 475 -181 479 -177
rect 495 -180 497 -176
rect 470 -182 479 -181
rect 477 -185 479 -182
rect 487 -185 489 -180
rect 495 -182 499 -180
rect 497 -185 499 -182
rect 504 -185 506 -176
rect 545 -180 547 -172
rect 561 -176 563 -172
rect 575 -175 576 -171
rect 580 -175 581 -171
rect 575 -176 581 -175
rect 585 -171 591 -170
rect 585 -175 586 -171
rect 590 -175 591 -171
rect 585 -176 591 -175
rect 615 -171 617 -168
rect 625 -171 627 -168
rect 615 -172 621 -171
rect 615 -176 616 -172
rect 620 -176 621 -172
rect 625 -174 629 -171
rect 554 -177 563 -176
rect 461 -192 463 -189
rect 461 -194 466 -192
rect 252 -204 254 -199
rect 259 -204 261 -199
rect 219 -206 244 -204
rect 298 -204 300 -199
rect 305 -204 307 -199
rect 395 -202 397 -197
rect 402 -202 404 -197
rect 464 -202 466 -194
rect 477 -198 479 -194
rect 487 -202 489 -194
rect 554 -181 555 -177
rect 559 -181 563 -177
rect 579 -180 581 -176
rect 554 -182 563 -181
rect 561 -185 563 -182
rect 571 -185 573 -180
rect 579 -182 583 -180
rect 581 -185 583 -182
rect 588 -185 590 -176
rect 615 -177 621 -176
rect 615 -185 617 -177
rect 545 -192 547 -189
rect 545 -194 550 -192
rect 497 -202 499 -197
rect 504 -202 506 -197
rect 464 -204 489 -202
rect 548 -202 550 -194
rect 561 -198 563 -194
rect 571 -202 573 -194
rect 627 -188 629 -174
rect 635 -179 637 -168
rect 710 -169 716 -168
rect 710 -173 711 -169
rect 715 -173 716 -169
rect 720 -171 724 -168
rect 710 -174 716 -173
rect 634 -180 640 -179
rect 634 -184 635 -180
rect 639 -184 640 -180
rect 710 -182 712 -174
rect 634 -185 640 -184
rect 634 -188 636 -185
rect 722 -185 724 -171
rect 730 -176 732 -165
rect 785 -167 787 -158
rect 832 -137 834 -133
rect 880 -137 882 -133
rect 812 -146 814 -142
rect 822 -146 824 -142
rect 865 -153 871 -152
rect 865 -157 866 -153
rect 870 -157 871 -153
rect 865 -158 871 -157
rect 796 -167 798 -164
rect 812 -167 814 -164
rect 822 -167 824 -164
rect 832 -167 834 -164
rect 785 -169 798 -167
rect 804 -169 814 -167
rect 818 -168 824 -167
rect 729 -177 735 -176
rect 788 -177 790 -169
rect 804 -173 806 -169
rect 818 -172 819 -168
rect 823 -172 824 -168
rect 818 -173 824 -172
rect 828 -168 834 -167
rect 828 -172 829 -168
rect 833 -172 834 -168
rect 869 -167 871 -158
rect 916 -137 918 -133
rect 896 -146 898 -142
rect 906 -146 908 -142
rect 1139 -139 1141 -136
rect 1178 -139 1180 -136
rect 1199 -139 1201 -136
rect 1232 -139 1234 -136
rect 1253 -139 1255 -136
rect 1288 -139 1290 -136
rect 1309 -139 1311 -136
rect 1342 -139 1344 -136
rect 1363 -139 1365 -136
rect 1694 -123 1700 -122
rect 1694 -125 1695 -123
rect 1668 -127 1673 -125
rect 1683 -127 1695 -125
rect 1699 -126 1700 -123
rect 1699 -127 1703 -126
rect 1694 -128 1703 -127
rect 1712 -128 1717 -126
rect 1662 -132 1668 -131
rect 1662 -136 1663 -132
rect 1667 -135 1668 -132
rect 1686 -135 1703 -133
rect 1712 -135 1717 -133
rect 1667 -136 1673 -135
rect 1662 -137 1673 -136
rect 1683 -137 1689 -135
rect 952 -145 958 -144
rect 942 -153 944 -148
rect 952 -149 953 -145
rect 957 -149 958 -145
rect 952 -150 958 -149
rect 880 -167 882 -164
rect 896 -167 898 -164
rect 906 -167 908 -164
rect 916 -167 918 -164
rect 952 -155 954 -150
rect 962 -155 964 -150
rect 1139 -160 1141 -142
rect 1178 -160 1180 -145
rect 1199 -160 1201 -145
rect 1232 -160 1234 -145
rect 1253 -160 1255 -145
rect 1288 -160 1290 -145
rect 1309 -160 1311 -145
rect 1342 -160 1344 -145
rect 1363 -160 1365 -145
rect 1686 -142 1692 -141
rect 1686 -145 1687 -142
rect 1666 -147 1671 -145
rect 1683 -146 1687 -145
rect 1691 -145 1692 -142
rect 1691 -146 1700 -145
rect 1683 -147 1700 -146
rect 1706 -147 1710 -145
rect 1580 -156 1584 -154
rect 1590 -155 1607 -154
rect 1590 -156 1599 -155
rect 1179 -164 1180 -160
rect 1200 -164 1201 -160
rect 1233 -164 1234 -160
rect 1254 -164 1255 -160
rect 1289 -164 1290 -160
rect 1310 -164 1311 -160
rect 1343 -164 1344 -160
rect 1364 -164 1365 -160
rect 1598 -159 1599 -156
rect 1603 -156 1607 -155
rect 1619 -156 1624 -154
rect 1603 -159 1604 -156
rect 1598 -160 1604 -159
rect 869 -169 882 -167
rect 888 -169 898 -167
rect 902 -168 908 -167
rect 828 -173 834 -172
rect 797 -174 806 -173
rect 729 -181 730 -177
rect 734 -181 735 -177
rect 729 -182 735 -181
rect 729 -185 731 -182
rect 615 -195 617 -191
rect 710 -192 712 -188
rect 797 -178 798 -174
rect 802 -178 806 -174
rect 822 -177 824 -173
rect 797 -179 806 -178
rect 804 -182 806 -179
rect 814 -182 816 -177
rect 822 -179 826 -177
rect 824 -182 826 -179
rect 831 -182 833 -173
rect 872 -177 874 -169
rect 888 -173 890 -169
rect 902 -172 903 -168
rect 907 -172 908 -168
rect 902 -173 908 -172
rect 912 -168 918 -167
rect 912 -172 913 -168
rect 917 -172 918 -168
rect 912 -173 918 -172
rect 942 -168 944 -165
rect 952 -168 954 -165
rect 942 -169 948 -168
rect 942 -173 943 -169
rect 947 -173 948 -169
rect 952 -171 956 -168
rect 881 -174 890 -173
rect 788 -189 790 -186
rect 788 -191 793 -189
rect 581 -202 583 -197
rect 588 -202 590 -197
rect 548 -204 573 -202
rect 627 -202 629 -197
rect 634 -202 636 -197
rect 722 -199 724 -194
rect 729 -199 731 -194
rect 791 -199 793 -191
rect 804 -195 806 -191
rect 814 -199 816 -191
rect 881 -178 882 -174
rect 886 -178 890 -174
rect 906 -177 908 -173
rect 881 -179 890 -178
rect 888 -182 890 -179
rect 898 -182 900 -177
rect 906 -179 910 -177
rect 908 -182 910 -179
rect 915 -182 917 -173
rect 942 -174 948 -173
rect 942 -182 944 -174
rect 872 -189 874 -186
rect 872 -191 877 -189
rect 824 -199 826 -194
rect 831 -199 833 -194
rect 791 -201 816 -199
rect 875 -199 877 -191
rect 888 -195 890 -191
rect 898 -199 900 -191
rect 954 -185 956 -171
rect 962 -176 964 -165
rect 1139 -176 1141 -164
rect 1178 -176 1180 -164
rect 1199 -176 1201 -164
rect 1232 -176 1234 -164
rect 1253 -176 1255 -164
rect 1288 -176 1290 -164
rect 1309 -176 1311 -164
rect 1342 -176 1344 -164
rect 1363 -176 1365 -164
rect 1601 -166 1607 -164
rect 1617 -165 1628 -164
rect 1617 -166 1623 -165
rect 1573 -168 1578 -166
rect 1587 -168 1604 -166
rect 1622 -169 1623 -166
rect 1627 -169 1628 -165
rect 1622 -170 1628 -169
rect 1573 -175 1578 -173
rect 1587 -174 1596 -173
rect 1587 -175 1591 -174
rect 961 -177 967 -176
rect 961 -181 962 -177
rect 966 -181 967 -177
rect 961 -182 967 -181
rect 1590 -178 1591 -175
rect 1595 -176 1607 -174
rect 1617 -176 1622 -174
rect 1595 -178 1596 -176
rect 1590 -179 1596 -178
rect 961 -185 963 -182
rect 942 -192 944 -188
rect 1139 -188 1141 -182
rect 1178 -188 1180 -182
rect 1199 -188 1201 -182
rect 1232 -188 1234 -182
rect 1253 -188 1255 -182
rect 1288 -188 1290 -182
rect 1309 -188 1311 -182
rect 1342 -188 1344 -182
rect 1363 -188 1365 -182
rect 908 -199 910 -194
rect 915 -199 917 -194
rect 875 -201 900 -199
rect 954 -199 956 -194
rect 961 -199 963 -194
rect 147 -221 149 -217
rect 157 -221 159 -217
rect 167 -221 169 -217
rect 476 -219 478 -215
rect 486 -219 488 -215
rect 496 -219 498 -215
rect 803 -216 805 -212
rect 813 -216 815 -212
rect 823 -216 825 -212
rect 1061 -222 1063 -220
rect 147 -235 149 -227
rect 143 -236 149 -235
rect 157 -236 159 -227
rect 167 -236 169 -227
rect 476 -233 478 -225
rect 143 -240 144 -236
rect 148 -240 149 -236
rect 163 -237 169 -236
rect 143 -241 149 -240
rect 147 -254 149 -241
rect 157 -243 159 -240
rect 163 -241 164 -237
rect 168 -241 169 -237
rect 472 -234 478 -233
rect 486 -234 488 -225
rect 496 -234 498 -225
rect 803 -230 805 -222
rect 472 -238 473 -234
rect 477 -238 478 -234
rect 492 -235 498 -234
rect 472 -239 478 -238
rect 163 -242 169 -241
rect 153 -244 159 -243
rect 153 -248 154 -244
rect 158 -248 159 -244
rect 153 -249 159 -248
rect 154 -254 156 -249
rect 167 -251 169 -242
rect 476 -252 478 -239
rect 486 -241 488 -238
rect 492 -239 493 -235
rect 497 -239 498 -235
rect 799 -231 805 -230
rect 813 -231 815 -222
rect 823 -231 825 -222
rect 1133 -222 1135 -216
rect 1172 -222 1174 -216
rect 1193 -222 1195 -216
rect 1226 -222 1228 -216
rect 1247 -222 1249 -216
rect 1282 -222 1284 -216
rect 1303 -222 1305 -216
rect 1336 -222 1338 -216
rect 1357 -222 1359 -216
rect 799 -235 800 -231
rect 804 -235 805 -231
rect 819 -232 825 -231
rect 799 -236 805 -235
rect 492 -240 498 -239
rect 482 -242 488 -241
rect 482 -246 483 -242
rect 487 -246 488 -242
rect 482 -247 488 -246
rect 483 -252 485 -247
rect 496 -249 498 -240
rect 803 -249 805 -236
rect 813 -238 815 -235
rect 819 -236 820 -232
rect 824 -236 825 -232
rect 819 -237 825 -236
rect 809 -239 815 -238
rect 809 -243 810 -239
rect 814 -243 815 -239
rect 809 -244 815 -243
rect 810 -249 812 -244
rect 823 -246 825 -237
rect 1061 -239 1063 -228
rect 1133 -240 1135 -228
rect 1172 -240 1174 -228
rect 1193 -240 1195 -228
rect 1226 -240 1228 -228
rect 1247 -240 1249 -228
rect 1282 -240 1284 -228
rect 1303 -240 1305 -228
rect 1336 -240 1338 -228
rect 1357 -240 1359 -228
rect 167 -267 169 -263
rect 496 -265 498 -261
rect 823 -262 825 -258
rect 1061 -261 1063 -243
rect 1173 -244 1174 -240
rect 1194 -244 1195 -240
rect 1227 -244 1228 -240
rect 1248 -244 1249 -240
rect 1283 -244 1284 -240
rect 1304 -244 1305 -240
rect 1337 -244 1338 -240
rect 1358 -244 1359 -240
rect 147 -276 149 -272
rect 154 -276 156 -272
rect 476 -274 478 -270
rect 483 -274 485 -270
rect 803 -271 805 -267
rect 810 -271 812 -267
rect 1061 -267 1063 -264
rect 1133 -262 1135 -244
rect 1172 -259 1174 -244
rect 1193 -259 1195 -244
rect 1226 -259 1228 -244
rect 1247 -259 1249 -244
rect 1282 -259 1284 -244
rect 1303 -259 1305 -244
rect 1336 -259 1338 -244
rect 1357 -259 1359 -244
rect 1415 -248 1417 -243
rect 1427 -244 1429 -239
rect 1686 -247 1692 -246
rect 1686 -249 1687 -247
rect 1660 -251 1665 -249
rect 1675 -251 1687 -249
rect 1691 -250 1692 -247
rect 1691 -251 1695 -250
rect 1686 -252 1695 -251
rect 1704 -252 1709 -250
rect 1415 -261 1417 -258
rect 1427 -261 1429 -258
rect 1411 -262 1417 -261
rect 1133 -268 1135 -265
rect 1172 -268 1174 -265
rect 1193 -268 1195 -265
rect 1226 -268 1228 -265
rect 1247 -268 1249 -265
rect 1282 -268 1284 -265
rect 1303 -268 1305 -265
rect 1336 -268 1338 -265
rect 1357 -268 1359 -265
rect 1411 -266 1412 -262
rect 1416 -266 1417 -262
rect 1411 -267 1417 -266
rect 1423 -262 1429 -261
rect 1423 -266 1424 -262
rect 1428 -266 1429 -262
rect 1423 -267 1429 -266
rect 1415 -270 1417 -267
rect 1427 -270 1429 -267
rect 1654 -256 1660 -255
rect 1654 -260 1655 -256
rect 1659 -259 1660 -256
rect 1678 -259 1695 -257
rect 1704 -259 1709 -257
rect 1659 -260 1665 -259
rect 1654 -261 1665 -260
rect 1675 -261 1681 -259
rect 139 -288 141 -284
rect 63 -296 69 -295
rect 53 -304 55 -299
rect 63 -300 64 -296
rect 68 -300 69 -296
rect 63 -301 69 -300
rect 63 -306 65 -301
rect 73 -306 75 -301
rect 124 -304 130 -303
rect 124 -308 125 -304
rect 129 -308 130 -304
rect 124 -309 130 -308
rect 53 -319 55 -316
rect 63 -319 65 -316
rect 53 -320 59 -319
rect 53 -324 54 -320
rect 58 -324 59 -320
rect 63 -322 67 -319
rect 53 -325 59 -324
rect 53 -333 55 -325
rect 65 -336 67 -322
rect 73 -327 75 -316
rect 128 -318 130 -309
rect 175 -288 177 -284
rect 223 -288 225 -284
rect 155 -297 157 -293
rect 165 -297 167 -293
rect 208 -304 214 -303
rect 208 -308 209 -304
rect 213 -308 214 -304
rect 208 -309 214 -308
rect 139 -318 141 -315
rect 155 -318 157 -315
rect 165 -318 167 -315
rect 175 -318 177 -315
rect 128 -320 141 -318
rect 147 -320 157 -318
rect 161 -319 167 -318
rect 72 -328 78 -327
rect 131 -328 133 -320
rect 147 -324 149 -320
rect 161 -323 162 -319
rect 166 -323 167 -319
rect 161 -324 167 -323
rect 171 -319 177 -318
rect 171 -323 172 -319
rect 176 -323 177 -319
rect 212 -318 214 -309
rect 259 -288 261 -284
rect 239 -297 241 -293
rect 249 -297 251 -293
rect 468 -286 470 -282
rect 392 -294 398 -293
rect 295 -296 301 -295
rect 285 -304 287 -299
rect 295 -300 296 -296
rect 300 -300 301 -296
rect 295 -301 301 -300
rect 223 -318 225 -315
rect 239 -318 241 -315
rect 249 -318 251 -315
rect 259 -318 261 -315
rect 295 -306 297 -301
rect 305 -306 307 -301
rect 382 -302 384 -297
rect 392 -298 393 -294
rect 397 -298 398 -294
rect 392 -299 398 -298
rect 392 -304 394 -299
rect 402 -304 404 -299
rect 453 -302 459 -301
rect 453 -306 454 -302
rect 458 -306 459 -302
rect 453 -307 459 -306
rect 212 -320 225 -318
rect 231 -320 241 -318
rect 245 -319 251 -318
rect 171 -324 177 -323
rect 140 -325 149 -324
rect 72 -332 73 -328
rect 77 -332 78 -328
rect 72 -333 78 -332
rect 72 -336 74 -333
rect 53 -343 55 -339
rect 140 -329 141 -325
rect 145 -329 149 -325
rect 165 -328 167 -324
rect 140 -330 149 -329
rect 147 -333 149 -330
rect 157 -333 159 -328
rect 165 -330 169 -328
rect 167 -333 169 -330
rect 174 -333 176 -324
rect 215 -328 217 -320
rect 231 -324 233 -320
rect 245 -323 246 -319
rect 250 -323 251 -319
rect 245 -324 251 -323
rect 255 -319 261 -318
rect 255 -323 256 -319
rect 260 -323 261 -319
rect 255 -324 261 -323
rect 285 -319 287 -316
rect 295 -319 297 -316
rect 285 -320 291 -319
rect 285 -324 286 -320
rect 290 -324 291 -320
rect 295 -322 299 -319
rect 224 -325 233 -324
rect 131 -340 133 -337
rect 131 -342 136 -340
rect 65 -350 67 -345
rect 72 -350 74 -345
rect 134 -350 136 -342
rect 147 -346 149 -342
rect 157 -350 159 -342
rect 224 -329 225 -325
rect 229 -329 233 -325
rect 249 -328 251 -324
rect 224 -330 233 -329
rect 231 -333 233 -330
rect 241 -333 243 -328
rect 249 -330 253 -328
rect 251 -333 253 -330
rect 258 -333 260 -324
rect 285 -325 291 -324
rect 285 -333 287 -325
rect 215 -340 217 -337
rect 215 -342 220 -340
rect 167 -350 169 -345
rect 174 -350 176 -345
rect 134 -352 159 -350
rect 218 -350 220 -342
rect 231 -346 233 -342
rect 241 -350 243 -342
rect 297 -336 299 -322
rect 305 -327 307 -316
rect 382 -317 384 -314
rect 392 -317 394 -314
rect 382 -318 388 -317
rect 382 -322 383 -318
rect 387 -322 388 -318
rect 392 -320 396 -317
rect 382 -323 388 -322
rect 304 -328 310 -327
rect 304 -332 305 -328
rect 309 -332 310 -328
rect 382 -331 384 -323
rect 304 -333 310 -332
rect 304 -336 306 -333
rect 285 -343 287 -339
rect 394 -334 396 -320
rect 402 -325 404 -314
rect 457 -316 459 -307
rect 504 -286 506 -282
rect 552 -286 554 -282
rect 484 -295 486 -291
rect 494 -295 496 -291
rect 537 -302 543 -301
rect 537 -306 538 -302
rect 542 -306 543 -302
rect 537 -307 543 -306
rect 468 -316 470 -313
rect 484 -316 486 -313
rect 494 -316 496 -313
rect 504 -316 506 -313
rect 457 -318 470 -316
rect 476 -318 486 -316
rect 490 -317 496 -316
rect 401 -326 407 -325
rect 460 -326 462 -318
rect 476 -322 478 -318
rect 490 -321 491 -317
rect 495 -321 496 -317
rect 490 -322 496 -321
rect 500 -317 506 -316
rect 500 -321 501 -317
rect 505 -321 506 -317
rect 541 -316 543 -307
rect 588 -286 590 -282
rect 568 -295 570 -291
rect 578 -295 580 -291
rect 795 -283 797 -279
rect 719 -291 725 -290
rect 624 -294 630 -293
rect 614 -302 616 -297
rect 624 -298 625 -294
rect 629 -298 630 -294
rect 624 -299 630 -298
rect 709 -299 711 -294
rect 719 -295 720 -291
rect 724 -295 725 -291
rect 719 -296 725 -295
rect 552 -316 554 -313
rect 568 -316 570 -313
rect 578 -316 580 -313
rect 588 -316 590 -313
rect 624 -304 626 -299
rect 634 -304 636 -299
rect 719 -301 721 -296
rect 729 -301 731 -296
rect 780 -299 786 -298
rect 780 -303 781 -299
rect 785 -303 786 -299
rect 780 -304 786 -303
rect 709 -314 711 -311
rect 719 -314 721 -311
rect 541 -318 554 -316
rect 560 -318 570 -316
rect 574 -317 580 -316
rect 500 -322 506 -321
rect 469 -323 478 -322
rect 401 -330 402 -326
rect 406 -330 407 -326
rect 401 -331 407 -330
rect 401 -334 403 -331
rect 382 -341 384 -337
rect 469 -327 470 -323
rect 474 -327 478 -323
rect 494 -326 496 -322
rect 469 -328 478 -327
rect 476 -331 478 -328
rect 486 -331 488 -326
rect 494 -328 498 -326
rect 496 -331 498 -328
rect 503 -331 505 -322
rect 544 -326 546 -318
rect 560 -322 562 -318
rect 574 -321 575 -317
rect 579 -321 580 -317
rect 574 -322 580 -321
rect 584 -317 590 -316
rect 584 -321 585 -317
rect 589 -321 590 -317
rect 584 -322 590 -321
rect 614 -317 616 -314
rect 624 -317 626 -314
rect 614 -318 620 -317
rect 614 -322 615 -318
rect 619 -322 620 -318
rect 624 -320 628 -317
rect 553 -323 562 -322
rect 460 -338 462 -335
rect 460 -340 465 -338
rect 251 -350 253 -345
rect 258 -350 260 -345
rect 218 -352 243 -350
rect 297 -350 299 -345
rect 304 -350 306 -345
rect 394 -348 396 -343
rect 401 -348 403 -343
rect 463 -348 465 -340
rect 476 -344 478 -340
rect 486 -348 488 -340
rect 553 -327 554 -323
rect 558 -327 562 -323
rect 578 -326 580 -322
rect 553 -328 562 -327
rect 560 -331 562 -328
rect 570 -331 572 -326
rect 578 -328 582 -326
rect 580 -331 582 -328
rect 587 -331 589 -322
rect 614 -323 620 -322
rect 614 -331 616 -323
rect 544 -338 546 -335
rect 544 -340 549 -338
rect 496 -348 498 -343
rect 503 -348 505 -343
rect 463 -350 488 -348
rect 547 -348 549 -340
rect 560 -344 562 -340
rect 570 -348 572 -340
rect 626 -334 628 -320
rect 634 -325 636 -314
rect 709 -315 715 -314
rect 709 -319 710 -315
rect 714 -319 715 -315
rect 719 -317 723 -314
rect 709 -320 715 -319
rect 633 -326 639 -325
rect 633 -330 634 -326
rect 638 -330 639 -326
rect 709 -328 711 -320
rect 633 -331 639 -330
rect 633 -334 635 -331
rect 721 -331 723 -317
rect 729 -322 731 -311
rect 784 -313 786 -304
rect 831 -283 833 -279
rect 879 -283 881 -279
rect 811 -292 813 -288
rect 821 -292 823 -288
rect 864 -299 870 -298
rect 864 -303 865 -299
rect 869 -303 870 -299
rect 864 -304 870 -303
rect 795 -313 797 -310
rect 811 -313 813 -310
rect 821 -313 823 -310
rect 831 -313 833 -310
rect 784 -315 797 -313
rect 803 -315 813 -313
rect 817 -314 823 -313
rect 728 -323 734 -322
rect 787 -323 789 -315
rect 803 -319 805 -315
rect 817 -318 818 -314
rect 822 -318 823 -314
rect 817 -319 823 -318
rect 827 -314 833 -313
rect 827 -318 828 -314
rect 832 -318 833 -314
rect 868 -313 870 -304
rect 915 -283 917 -279
rect 895 -292 897 -288
rect 905 -292 907 -288
rect 1137 -284 1139 -281
rect 1176 -284 1178 -281
rect 1197 -284 1199 -281
rect 1230 -284 1232 -281
rect 1251 -284 1253 -281
rect 1286 -284 1288 -281
rect 1307 -284 1309 -281
rect 1340 -284 1342 -281
rect 1361 -284 1363 -281
rect 951 -291 957 -290
rect 941 -299 943 -294
rect 951 -295 952 -291
rect 956 -295 957 -291
rect 951 -296 957 -295
rect 879 -313 881 -310
rect 895 -313 897 -310
rect 905 -313 907 -310
rect 915 -313 917 -310
rect 951 -301 953 -296
rect 961 -301 963 -296
rect 1137 -305 1139 -287
rect 1176 -305 1178 -290
rect 1197 -305 1199 -290
rect 1230 -305 1232 -290
rect 1251 -305 1253 -290
rect 1286 -305 1288 -290
rect 1307 -305 1309 -290
rect 1340 -305 1342 -290
rect 1361 -305 1363 -290
rect 1415 -292 1417 -287
rect 1678 -266 1684 -265
rect 1678 -269 1679 -266
rect 1658 -271 1663 -269
rect 1675 -270 1679 -269
rect 1683 -269 1684 -266
rect 1683 -270 1692 -269
rect 1675 -271 1692 -270
rect 1698 -271 1702 -269
rect 1643 -297 1647 -295
rect 1674 -296 1683 -295
rect 1674 -297 1678 -296
rect 1427 -302 1429 -298
rect 1677 -300 1678 -297
rect 1682 -298 1692 -296
rect 1704 -298 1709 -296
rect 1682 -300 1683 -298
rect 1677 -301 1683 -300
rect 1687 -305 1692 -303
rect 1704 -305 1709 -303
rect 1177 -309 1178 -305
rect 1198 -309 1199 -305
rect 1231 -309 1232 -305
rect 1252 -309 1253 -305
rect 1287 -309 1288 -305
rect 1308 -309 1309 -305
rect 1341 -309 1342 -305
rect 1362 -309 1363 -305
rect 1652 -307 1656 -305
rect 1674 -306 1689 -305
rect 1674 -307 1678 -306
rect 868 -315 881 -313
rect 887 -315 897 -313
rect 901 -314 907 -313
rect 827 -319 833 -318
rect 796 -320 805 -319
rect 728 -327 729 -323
rect 733 -327 734 -323
rect 728 -328 734 -327
rect 728 -331 730 -328
rect 614 -341 616 -337
rect 709 -338 711 -334
rect 796 -324 797 -320
rect 801 -324 805 -320
rect 821 -323 823 -319
rect 796 -325 805 -324
rect 803 -328 805 -325
rect 813 -328 815 -323
rect 821 -325 825 -323
rect 823 -328 825 -325
rect 830 -328 832 -319
rect 871 -323 873 -315
rect 887 -319 889 -315
rect 901 -318 902 -314
rect 906 -318 907 -314
rect 901 -319 907 -318
rect 911 -314 917 -313
rect 911 -318 912 -314
rect 916 -318 917 -314
rect 911 -319 917 -318
rect 941 -314 943 -311
rect 951 -314 953 -311
rect 941 -315 947 -314
rect 941 -319 942 -315
rect 946 -319 947 -315
rect 951 -317 955 -314
rect 880 -320 889 -319
rect 787 -335 789 -332
rect 787 -337 792 -335
rect 580 -348 582 -343
rect 587 -348 589 -343
rect 547 -350 572 -348
rect 626 -348 628 -343
rect 633 -348 635 -343
rect 721 -345 723 -340
rect 728 -345 730 -340
rect 790 -345 792 -337
rect 803 -341 805 -337
rect 813 -345 815 -337
rect 880 -324 881 -320
rect 885 -324 889 -320
rect 905 -323 907 -319
rect 880 -325 889 -324
rect 887 -328 889 -325
rect 897 -328 899 -323
rect 905 -325 909 -323
rect 907 -328 909 -325
rect 914 -328 916 -319
rect 941 -320 947 -319
rect 941 -328 943 -320
rect 871 -335 873 -332
rect 871 -337 876 -335
rect 823 -345 825 -340
rect 830 -345 832 -340
rect 790 -347 815 -345
rect 874 -345 876 -337
rect 887 -341 889 -337
rect 897 -345 899 -337
rect 953 -331 955 -317
rect 961 -322 963 -311
rect 1137 -321 1139 -309
rect 1176 -321 1178 -309
rect 1197 -321 1199 -309
rect 1230 -321 1232 -309
rect 1251 -321 1253 -309
rect 1286 -321 1288 -309
rect 1307 -321 1309 -309
rect 1340 -321 1342 -309
rect 1361 -321 1363 -309
rect 1677 -310 1678 -307
rect 1682 -307 1689 -306
rect 1682 -310 1683 -307
rect 1677 -311 1683 -310
rect 1687 -315 1692 -313
rect 1701 -315 1711 -313
rect 1652 -317 1656 -315
rect 1674 -317 1679 -315
rect 960 -323 966 -322
rect 960 -327 961 -323
rect 965 -327 966 -323
rect 1677 -323 1679 -317
rect 1677 -325 1692 -323
rect 1701 -325 1705 -323
rect 960 -328 966 -327
rect 960 -331 962 -328
rect 941 -338 943 -334
rect 1137 -333 1139 -327
rect 1176 -333 1178 -327
rect 1197 -333 1199 -327
rect 1230 -333 1232 -327
rect 1251 -333 1253 -327
rect 1286 -333 1288 -327
rect 1307 -333 1309 -327
rect 1340 -333 1342 -327
rect 1361 -333 1363 -327
rect 1429 -331 1431 -327
rect 1683 -327 1689 -325
rect 1683 -331 1684 -327
rect 1688 -331 1689 -327
rect 907 -345 909 -340
rect 914 -345 916 -340
rect 874 -347 899 -345
rect 953 -345 955 -340
rect 960 -345 962 -340
rect 1417 -342 1419 -337
rect 146 -367 148 -363
rect 156 -367 158 -363
rect 166 -367 168 -363
rect 475 -365 477 -361
rect 485 -365 487 -361
rect 495 -365 497 -361
rect 802 -362 804 -358
rect 812 -362 814 -358
rect 822 -362 824 -358
rect 1062 -364 1064 -362
rect 146 -381 148 -373
rect 142 -382 148 -381
rect 156 -382 158 -373
rect 166 -382 168 -373
rect 475 -379 477 -371
rect 142 -386 143 -382
rect 147 -386 148 -382
rect 162 -383 168 -382
rect 142 -387 148 -386
rect 146 -400 148 -387
rect 156 -389 158 -386
rect 162 -387 163 -383
rect 167 -387 168 -383
rect 471 -380 477 -379
rect 485 -380 487 -371
rect 495 -380 497 -371
rect 802 -376 804 -368
rect 471 -384 472 -380
rect 476 -384 477 -380
rect 491 -381 497 -380
rect 471 -385 477 -384
rect 162 -388 168 -387
rect 152 -390 158 -389
rect 152 -394 153 -390
rect 157 -394 158 -390
rect 152 -395 158 -394
rect 153 -400 155 -395
rect 166 -397 168 -388
rect 475 -398 477 -385
rect 485 -387 487 -384
rect 491 -385 492 -381
rect 496 -385 497 -381
rect 798 -377 804 -376
rect 812 -377 814 -368
rect 822 -377 824 -368
rect 1134 -364 1136 -358
rect 1173 -364 1175 -358
rect 1194 -364 1196 -358
rect 1227 -364 1229 -358
rect 1248 -364 1250 -358
rect 1283 -364 1285 -358
rect 1304 -364 1306 -358
rect 1337 -364 1339 -358
rect 1358 -364 1360 -358
rect 1643 -333 1647 -331
rect 1674 -333 1679 -331
rect 1683 -332 1689 -331
rect 1677 -339 1679 -333
rect 1709 -336 1711 -315
rect 1699 -338 1711 -336
rect 1699 -339 1701 -338
rect 1677 -341 1687 -339
rect 1696 -341 1701 -339
rect 1677 -342 1679 -341
rect 1662 -343 1679 -342
rect 1662 -347 1663 -343
rect 1667 -344 1679 -343
rect 1667 -347 1668 -344
rect 1662 -348 1668 -347
rect 1417 -362 1419 -359
rect 1429 -362 1431 -359
rect 1413 -363 1419 -362
rect 1413 -367 1414 -363
rect 1418 -367 1419 -363
rect 1413 -368 1419 -367
rect 1425 -363 1431 -362
rect 1425 -367 1426 -363
rect 1430 -367 1431 -363
rect 1425 -368 1431 -367
rect 798 -381 799 -377
rect 803 -381 804 -377
rect 818 -378 824 -377
rect 798 -382 804 -381
rect 491 -386 497 -385
rect 481 -388 487 -387
rect 481 -392 482 -388
rect 486 -392 487 -388
rect 481 -393 487 -392
rect 482 -398 484 -393
rect 495 -395 497 -386
rect 802 -395 804 -382
rect 812 -384 814 -381
rect 818 -382 819 -378
rect 823 -382 824 -378
rect 1062 -381 1064 -370
rect 818 -383 824 -382
rect 808 -385 814 -384
rect 808 -389 809 -385
rect 813 -389 814 -385
rect 808 -390 814 -389
rect 809 -395 811 -390
rect 822 -392 824 -383
rect 1134 -382 1136 -370
rect 1173 -382 1175 -370
rect 1194 -382 1196 -370
rect 1227 -382 1229 -370
rect 1248 -382 1250 -370
rect 1283 -382 1285 -370
rect 1304 -382 1306 -370
rect 1337 -382 1339 -370
rect 1358 -382 1360 -370
rect 1417 -371 1419 -368
rect 1429 -371 1431 -368
rect 166 -413 168 -409
rect 495 -411 497 -407
rect 822 -408 824 -404
rect 1062 -403 1064 -385
rect 1174 -386 1175 -382
rect 1195 -386 1196 -382
rect 1228 -386 1229 -382
rect 1249 -386 1250 -382
rect 1284 -386 1285 -382
rect 1305 -386 1306 -382
rect 1338 -386 1339 -382
rect 1359 -386 1360 -382
rect 1417 -386 1419 -381
rect 1643 -381 1647 -379
rect 1674 -380 1683 -379
rect 1674 -381 1678 -380
rect 1062 -409 1064 -406
rect 1134 -404 1136 -386
rect 1173 -401 1175 -386
rect 1194 -401 1196 -386
rect 1227 -401 1229 -386
rect 1248 -401 1250 -386
rect 1283 -401 1285 -386
rect 1304 -401 1306 -386
rect 1337 -401 1339 -386
rect 1358 -401 1360 -386
rect 1429 -390 1431 -385
rect 1677 -384 1678 -381
rect 1682 -382 1692 -380
rect 1704 -382 1709 -380
rect 1682 -384 1683 -382
rect 1677 -385 1683 -384
rect 1687 -389 1692 -387
rect 1704 -389 1709 -387
rect 1652 -391 1656 -389
rect 1674 -390 1689 -389
rect 1674 -391 1678 -390
rect 1677 -394 1678 -391
rect 1682 -391 1689 -390
rect 1682 -394 1683 -391
rect 1677 -395 1683 -394
rect 1687 -399 1692 -397
rect 1701 -399 1711 -397
rect 1652 -401 1656 -399
rect 1674 -401 1679 -399
rect 1134 -410 1136 -407
rect 1173 -410 1175 -407
rect 1194 -410 1196 -407
rect 1227 -410 1229 -407
rect 1248 -410 1250 -407
rect 1283 -410 1285 -407
rect 1304 -410 1306 -407
rect 1337 -410 1339 -407
rect 1358 -410 1360 -407
rect 1677 -407 1679 -401
rect 1677 -409 1692 -407
rect 1701 -409 1705 -407
rect 146 -422 148 -418
rect 153 -422 155 -418
rect 475 -420 477 -416
rect 482 -420 484 -416
rect 802 -417 804 -413
rect 809 -417 811 -413
rect 1683 -411 1689 -409
rect 1683 -415 1684 -411
rect 1688 -415 1689 -411
rect 1643 -417 1647 -415
rect 1674 -417 1679 -415
rect 1683 -416 1689 -415
rect 1138 -426 1140 -423
rect 1177 -426 1179 -423
rect 1198 -426 1200 -423
rect 1231 -426 1233 -423
rect 1252 -426 1254 -423
rect 1287 -426 1289 -423
rect 1308 -426 1310 -423
rect 1341 -426 1343 -423
rect 1362 -426 1364 -423
rect 347 -445 349 -441
rect 357 -443 359 -438
rect 367 -443 369 -438
rect 440 -445 442 -441
rect 450 -443 452 -438
rect 460 -443 462 -438
rect 347 -467 349 -463
rect 357 -467 359 -456
rect 367 -459 369 -456
rect 367 -460 373 -459
rect 367 -464 368 -460
rect 372 -464 373 -460
rect 527 -445 529 -441
rect 537 -443 539 -438
rect 547 -443 549 -438
rect 367 -465 373 -464
rect 347 -468 353 -467
rect 347 -472 348 -468
rect 352 -472 353 -468
rect 347 -473 353 -472
rect 357 -468 363 -467
rect 357 -472 358 -468
rect 362 -472 363 -468
rect 357 -473 363 -472
rect 347 -478 349 -473
rect 360 -478 362 -473
rect 367 -478 369 -465
rect 440 -467 442 -463
rect 450 -467 452 -456
rect 460 -459 462 -456
rect 460 -460 466 -459
rect 460 -464 461 -460
rect 465 -464 466 -460
rect 1138 -447 1140 -429
rect 1419 -427 1421 -422
rect 1431 -423 1433 -418
rect 1177 -447 1179 -432
rect 1198 -447 1200 -432
rect 1231 -447 1233 -432
rect 1252 -447 1254 -432
rect 1287 -447 1289 -432
rect 1308 -447 1310 -432
rect 1341 -447 1343 -432
rect 1362 -447 1364 -432
rect 1677 -423 1679 -417
rect 1709 -420 1711 -399
rect 1722 -390 1726 -388
rect 1732 -389 1756 -388
rect 1732 -390 1742 -389
rect 1741 -393 1742 -390
rect 1746 -390 1756 -389
rect 1768 -390 1772 -388
rect 1746 -393 1747 -390
rect 1741 -394 1747 -393
rect 1722 -400 1726 -398
rect 1732 -400 1741 -398
rect 1745 -399 1754 -398
rect 1745 -400 1749 -399
rect 1748 -403 1749 -400
rect 1753 -401 1754 -399
rect 1753 -403 1759 -401
rect 1777 -403 1781 -401
rect 1748 -404 1754 -403
rect 1722 -410 1726 -408
rect 1732 -409 1759 -408
rect 1732 -410 1741 -409
rect 1740 -413 1741 -410
rect 1745 -410 1759 -409
rect 1777 -410 1781 -408
rect 1745 -413 1746 -410
rect 1740 -414 1746 -413
rect 1699 -422 1711 -420
rect 1699 -423 1701 -422
rect 1677 -425 1687 -423
rect 1696 -425 1701 -423
rect 1677 -426 1679 -425
rect 1662 -427 1679 -426
rect 1662 -431 1663 -427
rect 1667 -428 1679 -427
rect 1667 -431 1668 -428
rect 1662 -432 1668 -431
rect 1419 -440 1421 -437
rect 1431 -440 1433 -437
rect 1712 -438 1716 -436
rect 1729 -437 1751 -436
rect 1729 -438 1733 -437
rect 1415 -441 1421 -440
rect 1415 -445 1416 -441
rect 1420 -445 1421 -441
rect 1415 -446 1421 -445
rect 1427 -441 1433 -440
rect 1427 -445 1428 -441
rect 1432 -445 1433 -441
rect 1427 -446 1433 -445
rect 1732 -441 1733 -438
rect 1737 -438 1751 -437
rect 1776 -438 1780 -436
rect 1737 -441 1738 -438
rect 1732 -442 1738 -441
rect 1742 -443 1748 -442
rect 1742 -446 1743 -443
rect 1178 -451 1179 -447
rect 1199 -451 1200 -447
rect 1232 -451 1233 -447
rect 1253 -451 1254 -447
rect 1288 -451 1289 -447
rect 1309 -451 1310 -447
rect 1342 -451 1343 -447
rect 1363 -451 1364 -447
rect 1419 -449 1421 -446
rect 1431 -449 1433 -446
rect 1714 -448 1719 -446
rect 1729 -447 1743 -446
rect 1747 -447 1748 -443
rect 1729 -448 1748 -447
rect 460 -465 466 -464
rect 440 -468 446 -467
rect 440 -472 441 -468
rect 445 -472 446 -468
rect 440 -473 446 -472
rect 450 -468 456 -467
rect 450 -472 451 -468
rect 455 -472 456 -468
rect 450 -473 456 -472
rect 440 -478 442 -473
rect 453 -478 455 -473
rect 460 -478 462 -465
rect 527 -467 529 -463
rect 537 -467 539 -456
rect 547 -459 549 -456
rect 547 -460 553 -459
rect 547 -464 548 -460
rect 552 -464 553 -460
rect 1138 -463 1140 -451
rect 1177 -463 1179 -451
rect 1198 -463 1200 -451
rect 1231 -463 1233 -451
rect 1252 -463 1254 -451
rect 1287 -463 1289 -451
rect 1308 -463 1310 -451
rect 1341 -463 1343 -451
rect 1362 -463 1364 -451
rect 547 -465 553 -464
rect 527 -468 533 -467
rect 527 -472 528 -468
rect 532 -472 533 -468
rect 527 -473 533 -472
rect 537 -468 543 -467
rect 537 -472 538 -468
rect 542 -472 543 -468
rect 537 -473 543 -472
rect 527 -478 529 -473
rect 540 -478 542 -473
rect 547 -478 549 -465
rect 1138 -475 1140 -469
rect 1177 -475 1179 -469
rect 1198 -475 1200 -469
rect 1231 -475 1233 -469
rect 1252 -475 1254 -469
rect 1287 -475 1289 -469
rect 1308 -475 1310 -469
rect 1341 -475 1343 -469
rect 1362 -475 1364 -469
rect 1419 -471 1421 -466
rect 347 -491 349 -487
rect 360 -494 362 -489
rect 367 -494 369 -489
rect 440 -491 442 -487
rect 453 -494 455 -489
rect 460 -494 462 -489
rect 527 -491 529 -487
rect 1746 -449 1748 -448
rect 1746 -451 1751 -449
rect 1764 -451 1769 -449
rect 1717 -458 1722 -456
rect 1736 -457 1745 -456
rect 1736 -458 1740 -457
rect 1739 -461 1740 -458
rect 1744 -459 1745 -457
rect 1744 -461 1748 -459
rect 1773 -461 1778 -459
rect 1739 -462 1745 -461
rect 1717 -468 1722 -466
rect 1736 -468 1748 -466
rect 1773 -468 1778 -466
rect 1431 -481 1433 -477
rect 540 -494 542 -489
rect 547 -494 549 -489
rect 1686 -479 1692 -478
rect 1686 -481 1687 -479
rect 1660 -483 1665 -481
rect 1675 -483 1687 -481
rect 1691 -482 1692 -479
rect 1739 -476 1745 -468
rect 1691 -483 1695 -482
rect 1686 -484 1695 -483
rect 1704 -484 1709 -482
rect 1739 -480 1740 -476
rect 1744 -480 1745 -476
rect 1654 -488 1660 -487
rect 1654 -492 1655 -488
rect 1659 -491 1660 -488
rect 1739 -483 1745 -480
rect 1739 -486 1740 -483
rect 1712 -488 1716 -486
rect 1736 -487 1740 -486
rect 1744 -484 1745 -483
rect 1744 -486 1748 -484
rect 1776 -486 1780 -484
rect 1744 -487 1745 -486
rect 1736 -488 1745 -487
rect 1678 -491 1695 -489
rect 1704 -491 1709 -489
rect 1659 -492 1665 -491
rect 1654 -493 1665 -492
rect 1675 -493 1681 -491
rect 1739 -493 1745 -492
rect 1678 -498 1684 -497
rect 1678 -501 1679 -498
rect 1658 -503 1663 -501
rect 1675 -502 1679 -501
rect 1683 -501 1684 -498
rect 1712 -495 1716 -493
rect 1736 -495 1740 -493
rect 1739 -497 1740 -495
rect 1744 -494 1745 -493
rect 1744 -496 1748 -494
rect 1776 -496 1784 -494
rect 1744 -497 1745 -496
rect 1739 -498 1745 -497
rect 1683 -502 1692 -501
rect 1675 -503 1692 -502
rect 1698 -503 1702 -501
rect 1739 -503 1745 -502
rect 1739 -504 1740 -503
rect 1714 -506 1716 -504
rect 1730 -506 1740 -504
rect 1739 -507 1740 -506
rect 1744 -504 1745 -503
rect 1744 -506 1748 -504
rect 1776 -506 1780 -504
rect 1744 -507 1745 -506
rect 1739 -508 1745 -507
rect 1782 -529 1784 -496
rect 1771 -531 1784 -529
rect 1771 -568 1773 -531
<< ndiffusion >>
rect 1701 472 1707 473
rect 1701 468 1702 472
rect 1706 471 1707 472
rect 1706 468 1710 471
rect 1701 466 1710 468
rect 1701 459 1710 464
rect 1701 455 1710 457
rect 132 445 139 446
rect 132 441 134 445
rect 138 441 139 445
rect 132 436 139 441
rect 219 445 226 446
rect 219 441 221 445
rect 225 441 226 445
rect 114 435 121 436
rect 114 431 115 435
rect 119 431 121 435
rect 114 430 121 431
rect 116 425 121 430
rect 123 425 128 436
rect 130 434 139 436
rect 219 436 226 441
rect 312 445 319 446
rect 312 441 314 445
rect 318 441 319 445
rect 201 435 208 436
rect 130 425 141 434
rect 143 433 150 434
rect 143 429 145 433
rect 149 429 150 433
rect 201 431 202 435
rect 206 431 208 435
rect 201 430 208 431
rect 143 428 150 429
rect 143 425 148 428
rect 203 425 208 430
rect 210 425 215 436
rect 217 434 226 436
rect 312 436 319 441
rect 545 447 552 448
rect 545 443 546 447
rect 550 443 552 447
rect 294 435 301 436
rect 217 425 228 434
rect 230 433 237 434
rect 230 429 232 433
rect 236 429 237 433
rect 294 431 295 435
rect 299 431 301 435
rect 294 430 301 431
rect 230 428 237 429
rect 230 425 235 428
rect 296 425 301 430
rect 303 425 308 436
rect 310 434 319 436
rect 545 438 552 443
rect 638 447 645 448
rect 638 443 639 447
rect 643 443 645 447
rect 545 436 554 438
rect 534 435 541 436
rect 310 425 321 434
rect 323 433 330 434
rect 323 429 325 433
rect 329 429 330 433
rect 534 431 535 435
rect 539 431 541 435
rect 534 430 541 431
rect 323 428 330 429
rect 323 425 328 428
rect 536 427 541 430
rect 543 427 554 436
rect 556 427 561 438
rect 563 437 570 438
rect 563 433 565 437
rect 569 433 570 437
rect 638 438 645 443
rect 725 447 732 448
rect 725 443 726 447
rect 730 443 732 447
rect 1582 444 1588 445
rect 638 436 647 438
rect 563 432 570 433
rect 627 435 634 436
rect 563 427 568 432
rect 627 431 628 435
rect 632 431 634 435
rect 627 430 634 431
rect 629 427 634 430
rect 636 427 647 436
rect 649 427 654 438
rect 656 437 663 438
rect 656 433 658 437
rect 662 433 663 437
rect 725 438 732 443
rect 725 436 734 438
rect 656 432 663 433
rect 714 435 721 436
rect 656 427 661 432
rect 714 431 715 435
rect 719 431 721 435
rect 714 430 721 431
rect 716 427 721 430
rect 723 427 734 436
rect 736 427 741 438
rect 743 437 750 438
rect 743 433 745 437
rect 749 433 750 437
rect 743 432 750 433
rect 743 427 748 432
rect 1582 440 1583 444
rect 1587 440 1588 444
rect 1582 438 1588 440
rect 1698 454 1716 455
rect 1698 450 1711 454
rect 1715 450 1716 454
rect 1698 449 1716 450
rect 1698 447 1704 449
rect 1582 434 1588 436
rect 1570 433 1588 434
rect 1570 429 1571 433
rect 1575 429 1588 433
rect 1570 428 1588 429
rect 1698 443 1704 445
rect 1698 439 1699 443
rect 1703 439 1704 443
rect 1698 438 1704 439
rect 1576 426 1585 428
rect 1576 419 1585 424
rect 1576 415 1585 417
rect 1576 412 1580 415
rect 1031 392 1042 395
rect 1044 392 1061 395
rect 1579 411 1580 412
rect 1584 411 1585 415
rect 1579 410 1585 411
rect 1698 427 1716 428
rect 1698 423 1711 427
rect 1715 423 1716 427
rect 1698 422 1716 423
rect 1698 420 1710 422
rect 1698 413 1710 418
rect 1698 409 1710 411
rect 1698 405 1701 409
rect 1705 406 1710 409
rect 1705 405 1707 406
rect 1698 403 1707 405
rect 1143 396 1153 397
rect 1103 391 1114 394
rect 1116 391 1133 394
rect 1143 392 1145 396
rect 1149 392 1153 396
rect 1143 391 1153 392
rect 1155 391 1174 397
rect 1176 396 1184 397
rect 1176 392 1179 396
rect 1183 392 1184 396
rect 1176 391 1184 392
rect 1197 396 1207 397
rect 1197 392 1199 396
rect 1203 392 1207 396
rect 1197 391 1207 392
rect 1209 391 1228 397
rect 1230 396 1238 397
rect 1230 392 1233 396
rect 1237 392 1238 396
rect 1230 391 1238 392
rect 1253 396 1263 397
rect 1253 392 1255 396
rect 1259 392 1263 396
rect 1253 391 1263 392
rect 1265 391 1284 397
rect 1286 396 1294 397
rect 1286 392 1289 396
rect 1293 392 1294 396
rect 1286 391 1294 392
rect 1307 396 1317 397
rect 1307 392 1309 396
rect 1313 392 1317 396
rect 1307 391 1317 392
rect 1319 391 1338 397
rect 1340 396 1348 397
rect 1340 392 1343 396
rect 1347 392 1348 396
rect 1340 391 1348 392
rect 1698 399 1707 401
rect 1698 395 1699 399
rect 1703 395 1707 399
rect 1698 393 1707 395
rect 1698 387 1707 391
rect 1698 383 1702 387
rect 1706 383 1707 387
rect 1698 382 1707 383
rect 1693 377 1702 382
rect 36 318 43 319
rect 36 314 37 318
rect 41 314 43 318
rect 36 313 43 314
rect 45 316 53 319
rect 114 323 121 324
rect 114 319 115 323
rect 119 319 121 323
rect 114 318 121 319
rect 45 313 55 316
rect 47 307 55 313
rect 57 307 62 316
rect 64 315 71 316
rect 116 315 121 318
rect 123 319 128 324
rect 198 323 205 324
rect 198 319 199 323
rect 203 319 205 323
rect 123 315 137 319
rect 64 311 66 315
rect 70 311 71 315
rect 64 310 71 311
rect 128 311 129 315
rect 133 311 137 315
rect 128 310 137 311
rect 139 318 147 319
rect 139 314 141 318
rect 145 314 147 318
rect 139 310 147 314
rect 149 316 157 319
rect 149 312 151 316
rect 155 312 157 316
rect 149 310 157 312
rect 64 307 69 310
rect 47 306 53 307
rect 47 302 48 306
rect 52 302 53 306
rect 47 301 53 302
rect 152 307 157 310
rect 159 307 164 319
rect 166 307 174 319
rect 198 318 205 319
rect 200 315 205 318
rect 207 319 212 324
rect 207 315 221 319
rect 212 311 213 315
rect 217 311 221 315
rect 212 310 221 311
rect 223 318 231 319
rect 223 314 225 318
rect 229 314 231 318
rect 223 310 231 314
rect 233 316 241 319
rect 233 312 235 316
rect 239 312 241 316
rect 233 310 241 312
rect 168 306 174 307
rect 168 302 169 306
rect 173 302 174 306
rect 168 301 174 302
rect 236 307 241 310
rect 243 307 248 319
rect 250 307 258 319
rect 268 318 275 319
rect 268 314 269 318
rect 273 314 275 318
rect 268 313 275 314
rect 277 316 285 319
rect 365 320 372 321
rect 365 316 366 320
rect 370 316 372 320
rect 277 313 287 316
rect 279 307 287 313
rect 289 307 294 316
rect 296 315 303 316
rect 365 315 372 316
rect 374 318 382 321
rect 443 325 450 326
rect 443 321 444 325
rect 448 321 450 325
rect 443 320 450 321
rect 374 315 384 318
rect 296 311 298 315
rect 302 311 303 315
rect 296 310 303 311
rect 296 307 301 310
rect 376 309 384 315
rect 386 309 391 318
rect 393 317 400 318
rect 445 317 450 320
rect 452 321 457 326
rect 527 325 534 326
rect 527 321 528 325
rect 532 321 534 325
rect 452 317 466 321
rect 393 313 395 317
rect 399 313 400 317
rect 393 312 400 313
rect 457 313 458 317
rect 462 313 466 317
rect 457 312 466 313
rect 468 320 476 321
rect 468 316 470 320
rect 474 316 476 320
rect 468 312 476 316
rect 478 318 486 321
rect 478 314 480 318
rect 484 314 486 318
rect 478 312 486 314
rect 393 309 398 312
rect 252 306 258 307
rect 252 302 253 306
rect 257 302 258 306
rect 252 301 258 302
rect 279 306 285 307
rect 279 302 280 306
rect 284 302 285 306
rect 376 308 382 309
rect 376 304 377 308
rect 381 304 382 308
rect 376 303 382 304
rect 481 309 486 312
rect 488 309 493 321
rect 495 309 503 321
rect 527 320 534 321
rect 529 317 534 320
rect 536 321 541 326
rect 536 317 550 321
rect 541 313 542 317
rect 546 313 550 317
rect 541 312 550 313
rect 552 320 560 321
rect 552 316 554 320
rect 558 316 560 320
rect 552 312 560 316
rect 562 318 570 321
rect 562 314 564 318
rect 568 314 570 318
rect 562 312 570 314
rect 497 308 503 309
rect 497 304 498 308
rect 502 304 503 308
rect 497 303 503 304
rect 565 309 570 312
rect 572 309 577 321
rect 579 309 587 321
rect 597 320 604 321
rect 597 316 598 320
rect 602 316 604 320
rect 597 315 604 316
rect 606 318 614 321
rect 692 323 699 324
rect 692 319 693 323
rect 697 319 699 323
rect 692 318 699 319
rect 701 321 709 324
rect 1107 369 1118 372
rect 1120 369 1137 372
rect 1147 371 1157 372
rect 1147 367 1149 371
rect 1153 367 1157 371
rect 1147 366 1157 367
rect 1159 366 1178 372
rect 1180 371 1188 372
rect 1180 367 1183 371
rect 1187 367 1188 371
rect 1180 366 1188 367
rect 1201 371 1211 372
rect 1201 367 1203 371
rect 1207 367 1211 371
rect 1201 366 1211 367
rect 1213 366 1232 372
rect 1234 371 1242 372
rect 1234 367 1237 371
rect 1241 367 1242 371
rect 1234 366 1242 367
rect 1257 371 1267 372
rect 1257 367 1259 371
rect 1263 367 1267 371
rect 1257 366 1267 367
rect 1269 366 1288 372
rect 1290 371 1298 372
rect 1290 367 1293 371
rect 1297 367 1298 371
rect 1290 366 1298 367
rect 1311 371 1321 372
rect 1311 367 1313 371
rect 1317 367 1321 371
rect 1311 366 1321 367
rect 1323 366 1342 372
rect 1344 371 1352 372
rect 1344 367 1347 371
rect 1351 367 1352 371
rect 1693 373 1702 375
rect 1693 369 1694 373
rect 1698 370 1702 373
rect 1698 369 1699 370
rect 1693 368 1699 369
rect 1344 366 1352 367
rect 1587 366 1593 367
rect 1587 365 1588 366
rect 1584 362 1588 365
rect 1592 362 1593 366
rect 1584 360 1593 362
rect 770 328 777 329
rect 770 324 771 328
rect 775 324 777 328
rect 770 323 777 324
rect 701 318 711 321
rect 606 315 616 318
rect 608 309 616 315
rect 618 309 623 318
rect 625 317 632 318
rect 625 313 627 317
rect 631 313 632 317
rect 625 312 632 313
rect 703 312 711 318
rect 713 312 718 321
rect 720 320 727 321
rect 772 320 777 323
rect 779 324 784 329
rect 854 328 861 329
rect 854 324 855 328
rect 859 324 861 328
rect 779 320 793 324
rect 720 316 722 320
rect 726 316 727 320
rect 720 315 727 316
rect 784 316 785 320
rect 789 316 793 320
rect 784 315 793 316
rect 795 323 803 324
rect 795 319 797 323
rect 801 319 803 323
rect 795 315 803 319
rect 805 321 813 324
rect 805 317 807 321
rect 811 317 813 321
rect 805 315 813 317
rect 720 312 725 315
rect 625 309 630 312
rect 581 308 587 309
rect 581 304 582 308
rect 586 304 587 308
rect 581 303 587 304
rect 608 308 614 309
rect 608 304 609 308
rect 613 304 614 308
rect 703 311 709 312
rect 703 307 704 311
rect 708 307 709 311
rect 703 306 709 307
rect 808 312 813 315
rect 815 312 820 324
rect 822 312 830 324
rect 854 323 861 324
rect 856 320 861 323
rect 863 324 868 329
rect 863 320 877 324
rect 868 316 869 320
rect 873 316 877 320
rect 868 315 877 316
rect 879 323 887 324
rect 879 319 881 323
rect 885 319 887 323
rect 879 315 887 319
rect 889 321 897 324
rect 889 317 891 321
rect 895 317 897 321
rect 889 315 897 317
rect 824 311 830 312
rect 824 307 825 311
rect 829 307 830 311
rect 824 306 830 307
rect 892 312 897 315
rect 899 312 904 324
rect 906 312 914 324
rect 924 323 931 324
rect 924 319 925 323
rect 929 319 931 323
rect 924 318 931 319
rect 933 321 941 324
rect 1548 351 1554 352
rect 1548 347 1549 351
rect 1553 347 1554 351
rect 1548 345 1554 347
rect 1548 341 1554 343
rect 1548 337 1549 341
rect 1553 337 1554 341
rect 1548 335 1554 337
rect 1548 331 1554 333
rect 1548 327 1549 331
rect 1553 327 1554 331
rect 1548 325 1554 327
rect 933 318 943 321
rect 935 312 943 318
rect 945 312 950 321
rect 952 320 959 321
rect 952 316 954 320
rect 958 316 959 320
rect 1548 321 1554 323
rect 1548 317 1549 321
rect 1553 317 1554 321
rect 1584 353 1593 358
rect 1579 352 1588 353
rect 1579 348 1580 352
rect 1584 348 1588 352
rect 1579 344 1588 348
rect 1579 340 1588 342
rect 1579 336 1583 340
rect 1587 336 1588 340
rect 1579 334 1588 336
rect 1698 343 1716 344
rect 1698 339 1711 343
rect 1715 339 1716 343
rect 1698 338 1716 339
rect 1698 336 1710 338
rect 1579 330 1588 332
rect 1579 329 1581 330
rect 1576 326 1581 329
rect 1585 326 1588 330
rect 1576 324 1588 326
rect 1732 334 1738 335
rect 1698 329 1710 334
rect 1576 317 1588 322
rect 1548 316 1554 317
rect 952 315 959 316
rect 1698 325 1710 327
rect 1698 321 1701 325
rect 1705 322 1710 325
rect 1705 321 1707 322
rect 1698 319 1707 321
rect 952 312 957 315
rect 1576 313 1588 315
rect 1570 312 1588 313
rect 908 311 914 312
rect 908 307 909 311
rect 913 307 914 311
rect 908 306 914 307
rect 935 311 941 312
rect 935 307 936 311
rect 940 307 941 311
rect 1570 308 1571 312
rect 1575 308 1588 312
rect 935 306 941 307
rect 608 303 614 304
rect 279 301 285 302
rect 1570 307 1588 308
rect 1698 315 1707 317
rect 1698 311 1699 315
rect 1703 311 1707 315
rect 1698 309 1707 311
rect 785 289 792 290
rect 458 286 465 287
rect 129 284 136 285
rect 129 280 130 284
rect 134 280 136 284
rect 129 279 136 280
rect 138 284 146 285
rect 138 280 140 284
rect 144 280 146 284
rect 138 279 146 280
rect 148 284 156 285
rect 148 280 150 284
rect 154 280 156 284
rect 148 279 156 280
rect 158 284 165 285
rect 158 280 160 284
rect 164 280 165 284
rect 458 282 459 286
rect 463 282 465 286
rect 458 281 465 282
rect 467 286 475 287
rect 467 282 469 286
rect 473 282 475 286
rect 467 281 475 282
rect 477 286 485 287
rect 477 282 479 286
rect 483 282 485 286
rect 477 281 485 282
rect 487 286 494 287
rect 487 282 489 286
rect 493 282 494 286
rect 785 285 786 289
rect 790 285 792 289
rect 785 284 792 285
rect 794 289 802 290
rect 794 285 796 289
rect 800 285 802 289
rect 794 284 802 285
rect 804 289 812 290
rect 804 285 806 289
rect 810 285 812 289
rect 804 284 812 285
rect 814 289 821 290
rect 814 285 816 289
rect 820 285 821 289
rect 814 284 821 285
rect 487 281 494 282
rect 158 279 165 280
rect 1698 303 1707 307
rect 1698 299 1702 303
rect 1706 299 1707 303
rect 1698 298 1707 299
rect 1693 293 1702 298
rect 1732 330 1733 334
rect 1737 330 1738 334
rect 1732 328 1738 330
rect 1732 324 1738 326
rect 1732 320 1733 324
rect 1737 320 1738 324
rect 1732 318 1738 320
rect 1732 314 1738 316
rect 1732 310 1733 314
rect 1737 310 1738 314
rect 1732 308 1738 310
rect 1732 304 1738 306
rect 1732 300 1733 304
rect 1737 300 1738 304
rect 1732 299 1738 300
rect 1693 289 1702 291
rect 1693 285 1694 289
rect 1698 286 1702 289
rect 1698 285 1699 286
rect 1693 284 1699 285
rect 1587 282 1593 283
rect 1587 281 1588 282
rect 1584 278 1588 281
rect 1592 278 1593 282
rect 1584 276 1593 278
rect 1031 247 1042 250
rect 1044 247 1061 250
rect 1376 263 1383 264
rect 1376 259 1377 263
rect 1381 259 1383 263
rect 1376 258 1383 259
rect 1378 254 1383 258
rect 1385 255 1395 264
rect 1385 254 1388 255
rect 1143 251 1153 252
rect 1103 246 1114 249
rect 1116 246 1133 249
rect 1143 247 1145 251
rect 1149 247 1153 251
rect 1143 246 1153 247
rect 1155 246 1174 252
rect 1176 251 1184 252
rect 1176 247 1179 251
rect 1183 247 1184 251
rect 1176 246 1184 247
rect 1197 251 1207 252
rect 1197 247 1199 251
rect 1203 247 1207 251
rect 1197 246 1207 247
rect 1209 246 1228 252
rect 1230 251 1238 252
rect 1230 247 1233 251
rect 1237 247 1238 251
rect 1230 246 1238 247
rect 1253 251 1263 252
rect 1253 247 1255 251
rect 1259 247 1263 251
rect 1253 246 1263 247
rect 1265 246 1284 252
rect 1286 251 1294 252
rect 1286 247 1289 251
rect 1293 247 1294 251
rect 1286 246 1294 247
rect 1307 251 1317 252
rect 1307 247 1309 251
rect 1313 247 1317 251
rect 1307 246 1317 247
rect 1319 246 1338 252
rect 1340 251 1348 252
rect 1340 247 1343 251
rect 1347 247 1348 251
rect 1387 251 1388 254
rect 1392 251 1395 255
rect 1387 250 1395 251
rect 1397 263 1404 264
rect 1397 259 1399 263
rect 1403 259 1404 263
rect 1397 256 1404 259
rect 1397 252 1399 256
rect 1403 252 1404 256
rect 1397 250 1404 252
rect 1584 269 1593 274
rect 1579 268 1588 269
rect 1579 264 1580 268
rect 1584 264 1588 268
rect 1579 260 1588 264
rect 1579 256 1588 258
rect 1579 252 1583 256
rect 1587 252 1588 256
rect 1579 250 1588 252
rect 1340 246 1348 247
rect 1579 246 1588 248
rect 1579 245 1581 246
rect 1576 242 1581 245
rect 1585 242 1588 246
rect 1576 240 1588 242
rect 35 172 42 173
rect 35 168 36 172
rect 40 168 42 172
rect 35 167 42 168
rect 44 170 52 173
rect 113 177 120 178
rect 113 173 114 177
rect 118 173 120 177
rect 113 172 120 173
rect 44 167 54 170
rect 46 161 54 167
rect 56 161 61 170
rect 63 169 70 170
rect 115 169 120 172
rect 122 173 127 178
rect 197 177 204 178
rect 197 173 198 177
rect 202 173 204 177
rect 122 169 136 173
rect 63 165 65 169
rect 69 165 70 169
rect 63 164 70 165
rect 127 165 128 169
rect 132 165 136 169
rect 127 164 136 165
rect 138 172 146 173
rect 138 168 140 172
rect 144 168 146 172
rect 138 164 146 168
rect 148 170 156 173
rect 148 166 150 170
rect 154 166 156 170
rect 148 164 156 166
rect 63 161 68 164
rect 46 160 52 161
rect 46 156 47 160
rect 51 156 52 160
rect 46 155 52 156
rect 151 161 156 164
rect 158 161 163 173
rect 165 161 173 173
rect 197 172 204 173
rect 199 169 204 172
rect 206 173 211 178
rect 206 169 220 173
rect 211 165 212 169
rect 216 165 220 169
rect 211 164 220 165
rect 222 172 230 173
rect 222 168 224 172
rect 228 168 230 172
rect 222 164 230 168
rect 232 170 240 173
rect 232 166 234 170
rect 238 166 240 170
rect 232 164 240 166
rect 167 160 173 161
rect 167 156 168 160
rect 172 156 173 160
rect 167 155 173 156
rect 235 161 240 164
rect 242 161 247 173
rect 249 161 257 173
rect 267 172 274 173
rect 267 168 268 172
rect 272 168 274 172
rect 267 167 274 168
rect 276 170 284 173
rect 364 174 371 175
rect 364 170 365 174
rect 369 170 371 174
rect 276 167 286 170
rect 278 161 286 167
rect 288 161 293 170
rect 295 169 302 170
rect 364 169 371 170
rect 373 172 381 175
rect 442 179 449 180
rect 442 175 443 179
rect 447 175 449 179
rect 442 174 449 175
rect 373 169 383 172
rect 295 165 297 169
rect 301 165 302 169
rect 295 164 302 165
rect 295 161 300 164
rect 375 163 383 169
rect 385 163 390 172
rect 392 171 399 172
rect 444 171 449 174
rect 451 175 456 180
rect 526 179 533 180
rect 526 175 527 179
rect 531 175 533 179
rect 451 171 465 175
rect 392 167 394 171
rect 398 167 399 171
rect 392 166 399 167
rect 456 167 457 171
rect 461 167 465 171
rect 456 166 465 167
rect 467 174 475 175
rect 467 170 469 174
rect 473 170 475 174
rect 467 166 475 170
rect 477 172 485 175
rect 477 168 479 172
rect 483 168 485 172
rect 477 166 485 168
rect 392 163 397 166
rect 251 160 257 161
rect 251 156 252 160
rect 256 156 257 160
rect 251 155 257 156
rect 278 160 284 161
rect 278 156 279 160
rect 283 156 284 160
rect 375 162 381 163
rect 375 158 376 162
rect 380 158 381 162
rect 375 157 381 158
rect 480 163 485 166
rect 487 163 492 175
rect 494 163 502 175
rect 526 174 533 175
rect 528 171 533 174
rect 535 175 540 180
rect 535 171 549 175
rect 540 167 541 171
rect 545 167 549 171
rect 540 166 549 167
rect 551 174 559 175
rect 551 170 553 174
rect 557 170 559 174
rect 551 166 559 170
rect 561 172 569 175
rect 561 168 563 172
rect 567 168 569 172
rect 561 166 569 168
rect 496 162 502 163
rect 496 158 497 162
rect 501 158 502 162
rect 496 157 502 158
rect 564 163 569 166
rect 571 163 576 175
rect 578 163 586 175
rect 596 174 603 175
rect 596 170 597 174
rect 601 170 603 174
rect 596 169 603 170
rect 605 172 613 175
rect 691 177 698 178
rect 691 173 692 177
rect 696 173 698 177
rect 691 172 698 173
rect 700 175 708 178
rect 1107 224 1118 227
rect 1120 224 1137 227
rect 1147 226 1157 227
rect 1147 222 1149 226
rect 1153 222 1157 226
rect 1147 221 1157 222
rect 1159 221 1178 227
rect 1180 226 1188 227
rect 1180 222 1183 226
rect 1187 222 1188 226
rect 1180 221 1188 222
rect 1201 226 1211 227
rect 1201 222 1203 226
rect 1207 222 1211 226
rect 1201 221 1211 222
rect 1213 221 1232 227
rect 1234 226 1242 227
rect 1234 222 1237 226
rect 1241 222 1242 226
rect 1234 221 1242 222
rect 1257 226 1267 227
rect 1257 222 1259 226
rect 1263 222 1267 226
rect 1257 221 1267 222
rect 1269 221 1288 227
rect 1290 226 1298 227
rect 1290 222 1293 226
rect 1297 222 1298 226
rect 1290 221 1298 222
rect 1311 226 1321 227
rect 1311 222 1313 226
rect 1317 222 1321 226
rect 1311 221 1321 222
rect 1323 221 1342 227
rect 1344 226 1352 227
rect 1344 222 1347 226
rect 1351 222 1352 226
rect 1576 233 1588 238
rect 1576 229 1588 231
rect 1388 228 1396 229
rect 1388 225 1389 228
rect 1344 221 1352 222
rect 1379 221 1384 225
rect 1377 220 1384 221
rect 1377 216 1378 220
rect 1382 216 1384 220
rect 1377 215 1384 216
rect 1386 224 1389 225
rect 1393 224 1396 228
rect 1386 215 1396 224
rect 1398 227 1405 229
rect 1398 223 1400 227
rect 1404 223 1405 227
rect 1570 228 1588 229
rect 1570 224 1571 228
rect 1575 224 1588 228
rect 1570 223 1588 224
rect 1701 240 1707 241
rect 1701 236 1702 240
rect 1706 239 1707 240
rect 1706 236 1710 239
rect 1701 234 1710 236
rect 1398 220 1405 223
rect 1398 216 1400 220
rect 1404 216 1405 220
rect 1398 215 1405 216
rect 1701 227 1710 232
rect 1701 223 1710 225
rect 1582 212 1588 213
rect 1582 208 1583 212
rect 1587 208 1588 212
rect 1582 206 1588 208
rect 1698 222 1716 223
rect 1698 218 1711 222
rect 1715 218 1716 222
rect 1698 217 1716 218
rect 1698 215 1704 217
rect 769 182 776 183
rect 769 178 770 182
rect 774 178 776 182
rect 769 177 776 178
rect 700 172 710 175
rect 605 169 615 172
rect 607 163 615 169
rect 617 163 622 172
rect 624 171 631 172
rect 624 167 626 171
rect 630 167 631 171
rect 624 166 631 167
rect 702 166 710 172
rect 712 166 717 175
rect 719 174 726 175
rect 771 174 776 177
rect 778 178 783 183
rect 853 182 860 183
rect 853 178 854 182
rect 858 178 860 182
rect 778 174 792 178
rect 719 170 721 174
rect 725 170 726 174
rect 719 169 726 170
rect 783 170 784 174
rect 788 170 792 174
rect 783 169 792 170
rect 794 177 802 178
rect 794 173 796 177
rect 800 173 802 177
rect 794 169 802 173
rect 804 175 812 178
rect 804 171 806 175
rect 810 171 812 175
rect 804 169 812 171
rect 719 166 724 169
rect 624 163 629 166
rect 580 162 586 163
rect 580 158 581 162
rect 585 158 586 162
rect 580 157 586 158
rect 607 162 613 163
rect 607 158 608 162
rect 612 158 613 162
rect 702 165 708 166
rect 702 161 703 165
rect 707 161 708 165
rect 702 160 708 161
rect 807 166 812 169
rect 814 166 819 178
rect 821 166 829 178
rect 853 177 860 178
rect 855 174 860 177
rect 862 178 867 183
rect 862 174 876 178
rect 867 170 868 174
rect 872 170 876 174
rect 867 169 876 170
rect 878 177 886 178
rect 878 173 880 177
rect 884 173 886 177
rect 878 169 886 173
rect 888 175 896 178
rect 888 171 890 175
rect 894 171 896 175
rect 888 169 896 171
rect 823 165 829 166
rect 823 161 824 165
rect 828 161 829 165
rect 823 160 829 161
rect 891 166 896 169
rect 898 166 903 178
rect 905 166 913 178
rect 923 177 930 178
rect 923 173 924 177
rect 928 173 930 177
rect 923 172 930 173
rect 932 175 940 178
rect 932 172 942 175
rect 934 166 942 172
rect 944 166 949 175
rect 951 174 958 175
rect 951 170 953 174
rect 957 170 958 174
rect 1582 202 1588 204
rect 1570 201 1588 202
rect 1570 197 1571 201
rect 1575 197 1588 201
rect 1570 196 1588 197
rect 1698 211 1704 213
rect 1698 207 1699 211
rect 1703 207 1704 211
rect 1698 206 1704 207
rect 1576 194 1585 196
rect 1576 187 1585 192
rect 1576 183 1585 185
rect 1576 180 1580 183
rect 1579 179 1580 180
rect 1584 179 1585 183
rect 1579 178 1585 179
rect 951 169 958 170
rect 951 166 956 169
rect 907 165 913 166
rect 907 161 908 165
rect 912 161 913 165
rect 907 160 913 161
rect 934 165 940 166
rect 934 161 935 165
rect 939 161 940 165
rect 934 160 940 161
rect 607 157 613 158
rect 278 155 284 156
rect 784 143 791 144
rect 457 140 464 141
rect 128 138 135 139
rect 128 134 129 138
rect 133 134 135 138
rect 128 133 135 134
rect 137 138 145 139
rect 137 134 139 138
rect 143 134 145 138
rect 137 133 145 134
rect 147 138 155 139
rect 147 134 149 138
rect 153 134 155 138
rect 147 133 155 134
rect 157 138 164 139
rect 157 134 159 138
rect 163 134 164 138
rect 457 136 458 140
rect 462 136 464 140
rect 457 135 464 136
rect 466 140 474 141
rect 466 136 468 140
rect 472 136 474 140
rect 466 135 474 136
rect 476 140 484 141
rect 476 136 478 140
rect 482 136 484 140
rect 476 135 484 136
rect 486 140 493 141
rect 486 136 488 140
rect 492 136 493 140
rect 784 139 785 143
rect 789 139 791 143
rect 784 138 791 139
rect 793 143 801 144
rect 793 139 795 143
rect 799 139 801 143
rect 793 138 801 139
rect 803 143 811 144
rect 803 139 805 143
rect 809 139 811 143
rect 803 138 811 139
rect 813 143 820 144
rect 813 139 815 143
rect 819 139 820 143
rect 813 138 820 139
rect 486 135 493 136
rect 157 133 164 134
rect 1030 105 1041 108
rect 1043 105 1060 108
rect 1376 123 1383 124
rect 1376 119 1377 123
rect 1381 119 1383 123
rect 1376 118 1383 119
rect 1378 114 1383 118
rect 1385 115 1395 124
rect 1385 114 1388 115
rect 1142 109 1152 110
rect 1102 104 1113 107
rect 1115 104 1132 107
rect 1142 105 1144 109
rect 1148 105 1152 109
rect 1142 104 1152 105
rect 1154 104 1173 110
rect 1175 109 1183 110
rect 1175 105 1178 109
rect 1182 105 1183 109
rect 1175 104 1183 105
rect 1196 109 1206 110
rect 1196 105 1198 109
rect 1202 105 1206 109
rect 1196 104 1206 105
rect 1208 104 1227 110
rect 1229 109 1237 110
rect 1229 105 1232 109
rect 1236 105 1237 109
rect 1229 104 1237 105
rect 1252 109 1262 110
rect 1252 105 1254 109
rect 1258 105 1262 109
rect 1252 104 1262 105
rect 1264 104 1283 110
rect 1285 109 1293 110
rect 1285 105 1288 109
rect 1292 105 1293 109
rect 1285 104 1293 105
rect 1306 109 1316 110
rect 1306 105 1308 109
rect 1312 105 1316 109
rect 1306 104 1316 105
rect 1318 104 1337 110
rect 1339 109 1347 110
rect 1387 111 1388 114
rect 1392 111 1395 115
rect 1387 110 1395 111
rect 1397 123 1404 124
rect 1397 119 1399 123
rect 1403 119 1404 123
rect 1397 116 1404 119
rect 1397 112 1399 116
rect 1403 112 1404 116
rect 1397 110 1404 112
rect 1339 105 1342 109
rect 1346 105 1347 109
rect 1339 104 1347 105
rect 1703 112 1709 113
rect 1703 108 1704 112
rect 1708 111 1709 112
rect 1708 108 1712 111
rect 1703 106 1712 108
rect 1703 99 1712 104
rect 1703 95 1712 97
rect 1106 82 1117 85
rect 1119 82 1136 85
rect 1146 84 1156 85
rect 1146 80 1148 84
rect 1152 80 1156 84
rect 1146 79 1156 80
rect 1158 79 1177 85
rect 1179 84 1187 85
rect 1179 80 1182 84
rect 1186 80 1187 84
rect 1179 79 1187 80
rect 1200 84 1210 85
rect 1200 80 1202 84
rect 1206 80 1210 84
rect 1200 79 1210 80
rect 1212 79 1231 85
rect 1233 84 1241 85
rect 1233 80 1236 84
rect 1240 80 1241 84
rect 1233 79 1241 80
rect 1256 84 1266 85
rect 1256 80 1258 84
rect 1262 80 1266 84
rect 1256 79 1266 80
rect 1268 79 1287 85
rect 1289 84 1297 85
rect 1289 80 1292 84
rect 1296 80 1297 84
rect 1289 79 1297 80
rect 1310 84 1320 85
rect 1310 80 1312 84
rect 1316 80 1320 84
rect 1310 79 1320 80
rect 1322 79 1341 85
rect 1343 84 1351 85
rect 1584 84 1590 85
rect 1343 80 1346 84
rect 1350 80 1351 84
rect 1343 79 1351 80
rect 1584 80 1585 84
rect 1589 80 1590 84
rect 1584 78 1590 80
rect 1700 94 1718 95
rect 1700 90 1713 94
rect 1717 90 1718 94
rect 1700 89 1718 90
rect 1700 87 1706 89
rect 1584 74 1590 76
rect 1572 73 1590 74
rect 1572 69 1573 73
rect 1577 69 1590 73
rect 1572 68 1590 69
rect 1700 83 1706 85
rect 1700 79 1701 83
rect 1705 79 1706 83
rect 1700 78 1706 79
rect 1578 66 1587 68
rect 1578 59 1587 64
rect 1578 55 1587 57
rect 1578 52 1582 55
rect 1581 51 1582 52
rect 1586 51 1587 55
rect 1581 50 1587 51
rect 1700 67 1718 68
rect 1700 63 1713 67
rect 1717 63 1718 67
rect 1700 62 1718 63
rect 1700 60 1712 62
rect 1700 53 1712 58
rect 1700 49 1712 51
rect 1700 45 1703 49
rect 1707 46 1712 49
rect 1707 45 1709 46
rect 1700 43 1709 45
rect 1700 39 1709 41
rect 1700 35 1701 39
rect 1705 35 1709 39
rect 1700 33 1709 35
rect 331 25 336 28
rect 329 24 336 25
rect 329 20 330 24
rect 334 20 336 24
rect 329 19 336 20
rect 338 19 349 28
rect 340 17 349 19
rect 351 17 356 28
rect 358 23 363 28
rect 424 25 429 28
rect 422 24 429 25
rect 358 22 365 23
rect 358 18 360 22
rect 364 18 365 22
rect 422 20 423 24
rect 427 20 429 24
rect 422 19 429 20
rect 431 19 442 28
rect 358 17 365 18
rect 340 12 347 17
rect 433 17 442 19
rect 444 17 449 28
rect 451 23 456 28
rect 511 25 516 28
rect 509 24 516 25
rect 451 22 458 23
rect 451 18 453 22
rect 457 18 458 22
rect 509 20 510 24
rect 514 20 516 24
rect 509 19 516 20
rect 518 19 529 28
rect 451 17 458 18
rect 340 8 341 12
rect 345 8 347 12
rect 340 7 347 8
rect 433 12 440 17
rect 520 17 529 19
rect 531 17 536 28
rect 538 23 543 28
rect 1700 27 1709 31
rect 538 22 545 23
rect 538 18 540 22
rect 544 18 545 22
rect 538 17 545 18
rect 433 8 434 12
rect 438 8 440 12
rect 433 7 440 8
rect 520 12 527 17
rect 1700 23 1704 27
rect 1708 23 1709 27
rect 1700 22 1709 23
rect 1695 17 1704 22
rect 520 8 521 12
rect 525 8 527 12
rect 1695 13 1704 15
rect 1695 9 1696 13
rect 1700 10 1704 13
rect 1700 9 1701 10
rect 1695 8 1701 9
rect 520 7 527 8
rect 1589 6 1595 7
rect 1589 5 1590 6
rect 1586 2 1590 5
rect 1594 2 1595 6
rect 1586 0 1595 2
rect 1550 -9 1556 -8
rect 1550 -13 1551 -9
rect 1555 -13 1556 -9
rect 1550 -15 1556 -13
rect 1550 -19 1556 -17
rect 1550 -23 1551 -19
rect 1555 -23 1556 -19
rect 1550 -25 1556 -23
rect 1550 -29 1556 -27
rect 1550 -33 1551 -29
rect 1555 -33 1556 -29
rect 1550 -35 1556 -33
rect 1550 -39 1556 -37
rect 1550 -43 1551 -39
rect 1555 -43 1556 -39
rect 1586 -7 1595 -2
rect 1581 -8 1590 -7
rect 1581 -12 1582 -8
rect 1586 -12 1590 -8
rect 1581 -16 1590 -12
rect 1581 -20 1590 -18
rect 1581 -24 1585 -20
rect 1589 -24 1590 -20
rect 1581 -26 1590 -24
rect 1700 -17 1718 -16
rect 1700 -21 1713 -17
rect 1717 -21 1718 -17
rect 1700 -22 1718 -21
rect 1700 -24 1712 -22
rect 1581 -30 1590 -28
rect 1581 -31 1583 -30
rect 1578 -34 1583 -31
rect 1587 -34 1590 -30
rect 1578 -36 1590 -34
rect 1734 -26 1740 -25
rect 1700 -31 1712 -26
rect 1578 -43 1590 -38
rect 1550 -44 1556 -43
rect 1700 -35 1712 -33
rect 1700 -39 1703 -35
rect 1707 -38 1712 -35
rect 1707 -39 1709 -38
rect 1700 -41 1709 -39
rect 1578 -47 1590 -45
rect 1572 -48 1590 -47
rect 1572 -52 1573 -48
rect 1577 -52 1590 -48
rect 1572 -53 1590 -52
rect 1700 -45 1709 -43
rect 1700 -49 1701 -45
rect 1705 -49 1709 -45
rect 1700 -51 1709 -49
rect 143 -61 150 -60
rect 143 -65 145 -61
rect 149 -65 150 -61
rect 143 -70 150 -65
rect 230 -61 237 -60
rect 230 -65 232 -61
rect 236 -65 237 -61
rect 125 -71 132 -70
rect 125 -75 126 -71
rect 130 -75 132 -71
rect 125 -76 132 -75
rect 127 -81 132 -76
rect 134 -81 139 -70
rect 141 -72 150 -70
rect 230 -70 237 -65
rect 323 -61 330 -60
rect 323 -65 325 -61
rect 329 -65 330 -61
rect 212 -71 219 -70
rect 141 -81 152 -72
rect 154 -73 161 -72
rect 154 -77 156 -73
rect 160 -77 161 -73
rect 212 -75 213 -71
rect 217 -75 219 -71
rect 212 -76 219 -75
rect 154 -78 161 -77
rect 154 -81 159 -78
rect 214 -81 219 -76
rect 221 -81 226 -70
rect 228 -72 237 -70
rect 323 -70 330 -65
rect 556 -59 563 -58
rect 556 -63 557 -59
rect 561 -63 563 -59
rect 305 -71 312 -70
rect 228 -81 239 -72
rect 241 -73 248 -72
rect 241 -77 243 -73
rect 247 -77 248 -73
rect 305 -75 306 -71
rect 310 -75 312 -71
rect 305 -76 312 -75
rect 241 -78 248 -77
rect 241 -81 246 -78
rect 307 -81 312 -76
rect 314 -81 319 -70
rect 321 -72 330 -70
rect 556 -68 563 -63
rect 649 -59 656 -58
rect 649 -63 650 -59
rect 654 -63 656 -59
rect 556 -70 565 -68
rect 545 -71 552 -70
rect 321 -81 332 -72
rect 334 -73 341 -72
rect 334 -77 336 -73
rect 340 -77 341 -73
rect 545 -75 546 -71
rect 550 -75 552 -71
rect 545 -76 552 -75
rect 334 -78 341 -77
rect 334 -81 339 -78
rect 547 -79 552 -76
rect 554 -79 565 -70
rect 567 -79 572 -68
rect 574 -69 581 -68
rect 574 -73 576 -69
rect 580 -73 581 -69
rect 649 -68 656 -63
rect 736 -59 743 -58
rect 736 -63 737 -59
rect 741 -63 743 -59
rect 1700 -57 1709 -53
rect 649 -70 658 -68
rect 574 -74 581 -73
rect 638 -71 645 -70
rect 574 -79 579 -74
rect 638 -75 639 -71
rect 643 -75 645 -71
rect 638 -76 645 -75
rect 640 -79 645 -76
rect 647 -79 658 -70
rect 660 -79 665 -68
rect 667 -69 674 -68
rect 667 -73 669 -69
rect 673 -73 674 -69
rect 736 -68 743 -63
rect 1700 -61 1704 -57
rect 1708 -61 1709 -57
rect 1700 -62 1709 -61
rect 1695 -67 1704 -62
rect 1734 -30 1735 -26
rect 1739 -30 1740 -26
rect 1734 -32 1740 -30
rect 1734 -36 1740 -34
rect 1734 -40 1735 -36
rect 1739 -40 1740 -36
rect 1734 -42 1740 -40
rect 1734 -46 1740 -44
rect 1734 -50 1735 -46
rect 1739 -50 1740 -46
rect 1734 -52 1740 -50
rect 1734 -56 1740 -54
rect 1734 -60 1735 -56
rect 1739 -60 1740 -56
rect 1734 -61 1740 -60
rect 736 -70 745 -68
rect 667 -74 674 -73
rect 725 -71 732 -70
rect 667 -79 672 -74
rect 725 -75 726 -71
rect 730 -75 732 -71
rect 725 -76 732 -75
rect 727 -79 732 -76
rect 734 -79 745 -70
rect 747 -79 752 -68
rect 754 -69 761 -68
rect 754 -73 756 -69
rect 760 -73 761 -69
rect 754 -74 761 -73
rect 754 -79 759 -74
rect 1695 -71 1704 -69
rect 1695 -75 1696 -71
rect 1700 -74 1704 -71
rect 1700 -75 1701 -74
rect 1695 -76 1701 -75
rect 1589 -78 1595 -77
rect 1589 -79 1590 -78
rect 1586 -82 1590 -79
rect 1594 -82 1595 -78
rect 1586 -84 1595 -82
rect 1052 -119 1063 -116
rect 1065 -119 1082 -116
rect 1586 -91 1595 -86
rect 1581 -92 1590 -91
rect 1581 -96 1582 -92
rect 1586 -96 1590 -92
rect 1581 -100 1590 -96
rect 1581 -104 1590 -102
rect 1581 -108 1585 -104
rect 1589 -108 1590 -104
rect 1581 -110 1590 -108
rect 1581 -114 1590 -112
rect 1164 -115 1174 -114
rect 1124 -120 1135 -117
rect 1137 -120 1154 -117
rect 1164 -119 1166 -115
rect 1170 -119 1174 -115
rect 1164 -120 1174 -119
rect 1176 -120 1195 -114
rect 1197 -115 1205 -114
rect 1197 -119 1200 -115
rect 1204 -119 1205 -115
rect 1197 -120 1205 -119
rect 1218 -115 1228 -114
rect 1218 -119 1220 -115
rect 1224 -119 1228 -115
rect 1218 -120 1228 -119
rect 1230 -120 1249 -114
rect 1251 -115 1259 -114
rect 1251 -119 1254 -115
rect 1258 -119 1259 -115
rect 1251 -120 1259 -119
rect 1274 -115 1284 -114
rect 1274 -119 1276 -115
rect 1280 -119 1284 -115
rect 1274 -120 1284 -119
rect 1286 -120 1305 -114
rect 1307 -115 1315 -114
rect 1307 -119 1310 -115
rect 1314 -119 1315 -115
rect 1307 -120 1315 -119
rect 1328 -115 1338 -114
rect 1328 -119 1330 -115
rect 1334 -119 1338 -115
rect 1328 -120 1338 -119
rect 1340 -120 1359 -114
rect 1361 -115 1369 -114
rect 1581 -115 1583 -114
rect 1361 -119 1364 -115
rect 1368 -119 1369 -115
rect 1361 -120 1369 -119
rect 1578 -118 1583 -115
rect 1587 -118 1590 -114
rect 1578 -120 1590 -118
rect 1578 -127 1590 -122
rect 1578 -131 1590 -129
rect 1572 -132 1590 -131
rect 47 -188 54 -187
rect 47 -192 48 -188
rect 52 -192 54 -188
rect 47 -193 54 -192
rect 56 -190 64 -187
rect 125 -183 132 -182
rect 125 -187 126 -183
rect 130 -187 132 -183
rect 125 -188 132 -187
rect 56 -193 66 -190
rect 58 -199 66 -193
rect 68 -199 73 -190
rect 75 -191 82 -190
rect 127 -191 132 -188
rect 134 -187 139 -182
rect 209 -183 216 -182
rect 209 -187 210 -183
rect 214 -187 216 -183
rect 134 -191 148 -187
rect 75 -195 77 -191
rect 81 -195 82 -191
rect 75 -196 82 -195
rect 139 -195 140 -191
rect 144 -195 148 -191
rect 139 -196 148 -195
rect 150 -188 158 -187
rect 150 -192 152 -188
rect 156 -192 158 -188
rect 150 -196 158 -192
rect 160 -190 168 -187
rect 160 -194 162 -190
rect 166 -194 168 -190
rect 160 -196 168 -194
rect 75 -199 80 -196
rect 58 -200 64 -199
rect 58 -204 59 -200
rect 63 -204 64 -200
rect 58 -205 64 -204
rect 163 -199 168 -196
rect 170 -199 175 -187
rect 177 -199 185 -187
rect 209 -188 216 -187
rect 211 -191 216 -188
rect 218 -187 223 -182
rect 218 -191 232 -187
rect 223 -195 224 -191
rect 228 -195 232 -191
rect 223 -196 232 -195
rect 234 -188 242 -187
rect 234 -192 236 -188
rect 240 -192 242 -188
rect 234 -196 242 -192
rect 244 -190 252 -187
rect 244 -194 246 -190
rect 250 -194 252 -190
rect 244 -196 252 -194
rect 179 -200 185 -199
rect 179 -204 180 -200
rect 184 -204 185 -200
rect 179 -205 185 -204
rect 247 -199 252 -196
rect 254 -199 259 -187
rect 261 -199 269 -187
rect 279 -188 286 -187
rect 279 -192 280 -188
rect 284 -192 286 -188
rect 279 -193 286 -192
rect 288 -190 296 -187
rect 376 -186 383 -185
rect 376 -190 377 -186
rect 381 -190 383 -186
rect 288 -193 298 -190
rect 290 -199 298 -193
rect 300 -199 305 -190
rect 307 -191 314 -190
rect 376 -191 383 -190
rect 385 -188 393 -185
rect 454 -181 461 -180
rect 454 -185 455 -181
rect 459 -185 461 -181
rect 454 -186 461 -185
rect 385 -191 395 -188
rect 307 -195 309 -191
rect 313 -195 314 -191
rect 307 -196 314 -195
rect 307 -199 312 -196
rect 387 -197 395 -191
rect 397 -197 402 -188
rect 404 -189 411 -188
rect 456 -189 461 -186
rect 463 -185 468 -180
rect 538 -181 545 -180
rect 538 -185 539 -181
rect 543 -185 545 -181
rect 463 -189 477 -185
rect 404 -193 406 -189
rect 410 -193 411 -189
rect 404 -194 411 -193
rect 468 -193 469 -189
rect 473 -193 477 -189
rect 468 -194 477 -193
rect 479 -186 487 -185
rect 479 -190 481 -186
rect 485 -190 487 -186
rect 479 -194 487 -190
rect 489 -188 497 -185
rect 489 -192 491 -188
rect 495 -192 497 -188
rect 489 -194 497 -192
rect 404 -197 409 -194
rect 263 -200 269 -199
rect 263 -204 264 -200
rect 268 -204 269 -200
rect 263 -205 269 -204
rect 290 -200 296 -199
rect 290 -204 291 -200
rect 295 -204 296 -200
rect 387 -198 393 -197
rect 387 -202 388 -198
rect 392 -202 393 -198
rect 387 -203 393 -202
rect 492 -197 497 -194
rect 499 -197 504 -185
rect 506 -197 514 -185
rect 538 -186 545 -185
rect 540 -189 545 -186
rect 547 -185 552 -180
rect 547 -189 561 -185
rect 552 -193 553 -189
rect 557 -193 561 -189
rect 552 -194 561 -193
rect 563 -186 571 -185
rect 563 -190 565 -186
rect 569 -190 571 -186
rect 563 -194 571 -190
rect 573 -188 581 -185
rect 573 -192 575 -188
rect 579 -192 581 -188
rect 573 -194 581 -192
rect 508 -198 514 -197
rect 508 -202 509 -198
rect 513 -202 514 -198
rect 508 -203 514 -202
rect 576 -197 581 -194
rect 583 -197 588 -185
rect 590 -197 598 -185
rect 608 -186 615 -185
rect 608 -190 609 -186
rect 613 -190 615 -186
rect 608 -191 615 -190
rect 617 -188 625 -185
rect 703 -183 710 -182
rect 703 -187 704 -183
rect 708 -187 710 -183
rect 703 -188 710 -187
rect 712 -185 720 -182
rect 1572 -136 1573 -132
rect 1577 -136 1590 -132
rect 1572 -137 1590 -136
rect 1703 -120 1709 -119
rect 1703 -124 1704 -120
rect 1708 -121 1709 -120
rect 1708 -124 1712 -121
rect 1703 -126 1712 -124
rect 1703 -133 1712 -128
rect 1703 -137 1712 -135
rect 1128 -142 1139 -139
rect 1141 -142 1158 -139
rect 1168 -140 1178 -139
rect 1168 -144 1170 -140
rect 1174 -144 1178 -140
rect 1168 -145 1178 -144
rect 1180 -145 1199 -139
rect 1201 -140 1209 -139
rect 1201 -144 1204 -140
rect 1208 -144 1209 -140
rect 1201 -145 1209 -144
rect 1222 -140 1232 -139
rect 1222 -144 1224 -140
rect 1228 -144 1232 -140
rect 1222 -145 1232 -144
rect 1234 -145 1253 -139
rect 1255 -140 1263 -139
rect 1255 -144 1258 -140
rect 1262 -144 1263 -140
rect 1255 -145 1263 -144
rect 1278 -140 1288 -139
rect 1278 -144 1280 -140
rect 1284 -144 1288 -140
rect 1278 -145 1288 -144
rect 1290 -145 1309 -139
rect 1311 -140 1319 -139
rect 1311 -144 1314 -140
rect 1318 -144 1319 -140
rect 1311 -145 1319 -144
rect 1332 -140 1342 -139
rect 1332 -144 1334 -140
rect 1338 -144 1342 -140
rect 1332 -145 1342 -144
rect 1344 -145 1363 -139
rect 1365 -140 1373 -139
rect 1365 -144 1368 -140
rect 1372 -144 1373 -140
rect 1365 -145 1373 -144
rect 1584 -148 1590 -147
rect 1584 -152 1585 -148
rect 1589 -152 1590 -148
rect 1584 -154 1590 -152
rect 1700 -138 1718 -137
rect 1700 -142 1713 -138
rect 1717 -142 1718 -138
rect 1700 -143 1718 -142
rect 1700 -145 1706 -143
rect 1584 -158 1590 -156
rect 1572 -159 1590 -158
rect 1572 -163 1573 -159
rect 1577 -163 1590 -159
rect 1572 -164 1590 -163
rect 1700 -149 1706 -147
rect 1700 -153 1701 -149
rect 1705 -153 1706 -149
rect 1700 -154 1706 -153
rect 781 -178 788 -177
rect 781 -182 782 -178
rect 786 -182 788 -178
rect 781 -183 788 -182
rect 712 -188 722 -185
rect 617 -191 627 -188
rect 619 -197 627 -191
rect 629 -197 634 -188
rect 636 -189 643 -188
rect 636 -193 638 -189
rect 642 -193 643 -189
rect 636 -194 643 -193
rect 714 -194 722 -188
rect 724 -194 729 -185
rect 731 -186 738 -185
rect 783 -186 788 -183
rect 790 -182 795 -177
rect 865 -178 872 -177
rect 865 -182 866 -178
rect 870 -182 872 -178
rect 790 -186 804 -182
rect 731 -190 733 -186
rect 737 -190 738 -186
rect 731 -191 738 -190
rect 795 -190 796 -186
rect 800 -190 804 -186
rect 795 -191 804 -190
rect 806 -183 814 -182
rect 806 -187 808 -183
rect 812 -187 814 -183
rect 806 -191 814 -187
rect 816 -185 824 -182
rect 816 -189 818 -185
rect 822 -189 824 -185
rect 816 -191 824 -189
rect 731 -194 736 -191
rect 636 -197 641 -194
rect 592 -198 598 -197
rect 592 -202 593 -198
rect 597 -202 598 -198
rect 592 -203 598 -202
rect 619 -198 625 -197
rect 619 -202 620 -198
rect 624 -202 625 -198
rect 714 -195 720 -194
rect 714 -199 715 -195
rect 719 -199 720 -195
rect 714 -200 720 -199
rect 819 -194 824 -191
rect 826 -194 831 -182
rect 833 -194 841 -182
rect 865 -183 872 -182
rect 867 -186 872 -183
rect 874 -182 879 -177
rect 874 -186 888 -182
rect 879 -190 880 -186
rect 884 -190 888 -186
rect 879 -191 888 -190
rect 890 -183 898 -182
rect 890 -187 892 -183
rect 896 -187 898 -183
rect 890 -191 898 -187
rect 900 -185 908 -182
rect 900 -189 902 -185
rect 906 -189 908 -185
rect 900 -191 908 -189
rect 835 -195 841 -194
rect 835 -199 836 -195
rect 840 -199 841 -195
rect 835 -200 841 -199
rect 903 -194 908 -191
rect 910 -194 915 -182
rect 917 -194 925 -182
rect 935 -183 942 -182
rect 935 -187 936 -183
rect 940 -187 942 -183
rect 935 -188 942 -187
rect 944 -185 952 -182
rect 1578 -166 1587 -164
rect 1578 -173 1587 -168
rect 1578 -177 1587 -175
rect 1578 -180 1582 -177
rect 1581 -181 1582 -180
rect 1586 -181 1587 -177
rect 1581 -182 1587 -181
rect 944 -188 954 -185
rect 946 -194 954 -188
rect 956 -194 961 -185
rect 963 -186 970 -185
rect 963 -190 965 -186
rect 969 -190 970 -186
rect 963 -191 970 -190
rect 963 -194 968 -191
rect 919 -195 925 -194
rect 919 -199 920 -195
rect 924 -199 925 -195
rect 919 -200 925 -199
rect 946 -195 952 -194
rect 946 -199 947 -195
rect 951 -199 952 -195
rect 946 -200 952 -199
rect 619 -203 625 -202
rect 290 -205 296 -204
rect 796 -217 803 -216
rect 469 -220 476 -219
rect 140 -222 147 -221
rect 140 -226 141 -222
rect 145 -226 147 -222
rect 140 -227 147 -226
rect 149 -222 157 -221
rect 149 -226 151 -222
rect 155 -226 157 -222
rect 149 -227 157 -226
rect 159 -222 167 -221
rect 159 -226 161 -222
rect 165 -226 167 -222
rect 159 -227 167 -226
rect 169 -222 176 -221
rect 169 -226 171 -222
rect 175 -226 176 -222
rect 469 -224 470 -220
rect 474 -224 476 -220
rect 469 -225 476 -224
rect 478 -220 486 -219
rect 478 -224 480 -220
rect 484 -224 486 -220
rect 478 -225 486 -224
rect 488 -220 496 -219
rect 488 -224 490 -220
rect 494 -224 496 -220
rect 488 -225 496 -224
rect 498 -220 505 -219
rect 498 -224 500 -220
rect 504 -224 505 -220
rect 796 -221 797 -217
rect 801 -221 803 -217
rect 796 -222 803 -221
rect 805 -217 813 -216
rect 805 -221 807 -217
rect 811 -221 813 -217
rect 805 -222 813 -221
rect 815 -217 823 -216
rect 815 -221 817 -217
rect 821 -221 823 -217
rect 815 -222 823 -221
rect 825 -217 832 -216
rect 825 -221 827 -217
rect 831 -221 832 -217
rect 825 -222 832 -221
rect 498 -225 505 -224
rect 169 -227 176 -226
rect 1050 -264 1061 -261
rect 1063 -264 1080 -261
rect 1419 -245 1427 -244
rect 1419 -248 1420 -245
rect 1410 -252 1415 -248
rect 1408 -253 1415 -252
rect 1408 -257 1409 -253
rect 1413 -257 1415 -253
rect 1408 -258 1415 -257
rect 1417 -249 1420 -248
rect 1424 -249 1427 -245
rect 1417 -258 1427 -249
rect 1429 -246 1436 -244
rect 1429 -250 1431 -246
rect 1435 -250 1436 -246
rect 1429 -253 1436 -250
rect 1429 -257 1431 -253
rect 1435 -257 1436 -253
rect 1429 -258 1436 -257
rect 1695 -244 1701 -243
rect 1695 -248 1696 -244
rect 1700 -245 1701 -244
rect 1700 -248 1704 -245
rect 1695 -250 1704 -248
rect 1162 -260 1172 -259
rect 1122 -265 1133 -262
rect 1135 -265 1152 -262
rect 1162 -264 1164 -260
rect 1168 -264 1172 -260
rect 1162 -265 1172 -264
rect 1174 -265 1193 -259
rect 1195 -260 1203 -259
rect 1195 -264 1198 -260
rect 1202 -264 1203 -260
rect 1195 -265 1203 -264
rect 1216 -260 1226 -259
rect 1216 -264 1218 -260
rect 1222 -264 1226 -260
rect 1216 -265 1226 -264
rect 1228 -265 1247 -259
rect 1249 -260 1257 -259
rect 1249 -264 1252 -260
rect 1256 -264 1257 -260
rect 1249 -265 1257 -264
rect 1272 -260 1282 -259
rect 1272 -264 1274 -260
rect 1278 -264 1282 -260
rect 1272 -265 1282 -264
rect 1284 -265 1303 -259
rect 1305 -260 1313 -259
rect 1305 -264 1308 -260
rect 1312 -264 1313 -260
rect 1305 -265 1313 -264
rect 1326 -260 1336 -259
rect 1326 -264 1328 -260
rect 1332 -264 1336 -260
rect 1326 -265 1336 -264
rect 1338 -265 1357 -259
rect 1359 -260 1367 -259
rect 1359 -264 1362 -260
rect 1366 -264 1367 -260
rect 1359 -265 1367 -264
rect 1695 -257 1704 -252
rect 1695 -261 1704 -259
rect 46 -334 53 -333
rect 46 -338 47 -334
rect 51 -338 53 -334
rect 46 -339 53 -338
rect 55 -336 63 -333
rect 124 -329 131 -328
rect 124 -333 125 -329
rect 129 -333 131 -329
rect 124 -334 131 -333
rect 55 -339 65 -336
rect 57 -345 65 -339
rect 67 -345 72 -336
rect 74 -337 81 -336
rect 126 -337 131 -334
rect 133 -333 138 -328
rect 208 -329 215 -328
rect 208 -333 209 -329
rect 213 -333 215 -329
rect 133 -337 147 -333
rect 74 -341 76 -337
rect 80 -341 81 -337
rect 74 -342 81 -341
rect 138 -341 139 -337
rect 143 -341 147 -337
rect 138 -342 147 -341
rect 149 -334 157 -333
rect 149 -338 151 -334
rect 155 -338 157 -334
rect 149 -342 157 -338
rect 159 -336 167 -333
rect 159 -340 161 -336
rect 165 -340 167 -336
rect 159 -342 167 -340
rect 74 -345 79 -342
rect 57 -346 63 -345
rect 57 -350 58 -346
rect 62 -350 63 -346
rect 57 -351 63 -350
rect 162 -345 167 -342
rect 169 -345 174 -333
rect 176 -345 184 -333
rect 208 -334 215 -333
rect 210 -337 215 -334
rect 217 -333 222 -328
rect 217 -337 231 -333
rect 222 -341 223 -337
rect 227 -341 231 -337
rect 222 -342 231 -341
rect 233 -334 241 -333
rect 233 -338 235 -334
rect 239 -338 241 -334
rect 233 -342 241 -338
rect 243 -336 251 -333
rect 243 -340 245 -336
rect 249 -340 251 -336
rect 243 -342 251 -340
rect 178 -346 184 -345
rect 178 -350 179 -346
rect 183 -350 184 -346
rect 178 -351 184 -350
rect 246 -345 251 -342
rect 253 -345 258 -333
rect 260 -345 268 -333
rect 278 -334 285 -333
rect 278 -338 279 -334
rect 283 -338 285 -334
rect 278 -339 285 -338
rect 287 -336 295 -333
rect 375 -332 382 -331
rect 375 -336 376 -332
rect 380 -336 382 -332
rect 287 -339 297 -336
rect 289 -345 297 -339
rect 299 -345 304 -336
rect 306 -337 313 -336
rect 375 -337 382 -336
rect 384 -334 392 -331
rect 453 -327 460 -326
rect 453 -331 454 -327
rect 458 -331 460 -327
rect 453 -332 460 -331
rect 384 -337 394 -334
rect 306 -341 308 -337
rect 312 -341 313 -337
rect 306 -342 313 -341
rect 306 -345 311 -342
rect 386 -343 394 -337
rect 396 -343 401 -334
rect 403 -335 410 -334
rect 455 -335 460 -332
rect 462 -331 467 -326
rect 537 -327 544 -326
rect 537 -331 538 -327
rect 542 -331 544 -327
rect 462 -335 476 -331
rect 403 -339 405 -335
rect 409 -339 410 -335
rect 403 -340 410 -339
rect 467 -339 468 -335
rect 472 -339 476 -335
rect 467 -340 476 -339
rect 478 -332 486 -331
rect 478 -336 480 -332
rect 484 -336 486 -332
rect 478 -340 486 -336
rect 488 -334 496 -331
rect 488 -338 490 -334
rect 494 -338 496 -334
rect 488 -340 496 -338
rect 403 -343 408 -340
rect 262 -346 268 -345
rect 262 -350 263 -346
rect 267 -350 268 -346
rect 262 -351 268 -350
rect 289 -346 295 -345
rect 289 -350 290 -346
rect 294 -350 295 -346
rect 386 -344 392 -343
rect 386 -348 387 -344
rect 391 -348 392 -344
rect 386 -349 392 -348
rect 491 -343 496 -340
rect 498 -343 503 -331
rect 505 -343 513 -331
rect 537 -332 544 -331
rect 539 -335 544 -332
rect 546 -331 551 -326
rect 546 -335 560 -331
rect 551 -339 552 -335
rect 556 -339 560 -335
rect 551 -340 560 -339
rect 562 -332 570 -331
rect 562 -336 564 -332
rect 568 -336 570 -332
rect 562 -340 570 -336
rect 572 -334 580 -331
rect 572 -338 574 -334
rect 578 -338 580 -334
rect 572 -340 580 -338
rect 507 -344 513 -343
rect 507 -348 508 -344
rect 512 -348 513 -344
rect 507 -349 513 -348
rect 575 -343 580 -340
rect 582 -343 587 -331
rect 589 -343 597 -331
rect 607 -332 614 -331
rect 607 -336 608 -332
rect 612 -336 614 -332
rect 607 -337 614 -336
rect 616 -334 624 -331
rect 702 -329 709 -328
rect 702 -333 703 -329
rect 707 -333 709 -329
rect 702 -334 709 -333
rect 711 -331 719 -328
rect 1126 -287 1137 -284
rect 1139 -287 1156 -284
rect 1166 -285 1176 -284
rect 1166 -289 1168 -285
rect 1172 -289 1176 -285
rect 1166 -290 1176 -289
rect 1178 -290 1197 -284
rect 1199 -285 1207 -284
rect 1199 -289 1202 -285
rect 1206 -289 1207 -285
rect 1199 -290 1207 -289
rect 1220 -285 1230 -284
rect 1220 -289 1222 -285
rect 1226 -289 1230 -285
rect 1220 -290 1230 -289
rect 1232 -290 1251 -284
rect 1253 -285 1261 -284
rect 1253 -289 1256 -285
rect 1260 -289 1261 -285
rect 1253 -290 1261 -289
rect 1276 -285 1286 -284
rect 1276 -289 1278 -285
rect 1282 -289 1286 -285
rect 1276 -290 1286 -289
rect 1288 -290 1307 -284
rect 1309 -285 1317 -284
rect 1309 -289 1312 -285
rect 1316 -289 1317 -285
rect 1309 -290 1317 -289
rect 1330 -285 1340 -284
rect 1330 -289 1332 -285
rect 1336 -289 1340 -285
rect 1330 -290 1340 -289
rect 1342 -290 1361 -284
rect 1363 -285 1371 -284
rect 1363 -289 1366 -285
rect 1370 -289 1371 -285
rect 1363 -290 1371 -289
rect 1692 -262 1710 -261
rect 1692 -266 1705 -262
rect 1709 -266 1710 -262
rect 1692 -267 1710 -266
rect 1692 -269 1698 -267
rect 1692 -273 1698 -271
rect 1692 -277 1693 -273
rect 1697 -277 1698 -273
rect 1692 -278 1698 -277
rect 1692 -289 1710 -288
rect 1692 -293 1705 -289
rect 1709 -293 1710 -289
rect 1692 -294 1710 -293
rect 1692 -296 1704 -294
rect 1692 -303 1704 -298
rect 780 -324 787 -323
rect 780 -328 781 -324
rect 785 -328 787 -324
rect 780 -329 787 -328
rect 711 -334 721 -331
rect 616 -337 626 -334
rect 618 -343 626 -337
rect 628 -343 633 -334
rect 635 -335 642 -334
rect 635 -339 637 -335
rect 641 -339 642 -335
rect 635 -340 642 -339
rect 713 -340 721 -334
rect 723 -340 728 -331
rect 730 -332 737 -331
rect 782 -332 787 -329
rect 789 -328 794 -323
rect 864 -324 871 -323
rect 864 -328 865 -324
rect 869 -328 871 -324
rect 789 -332 803 -328
rect 730 -336 732 -332
rect 736 -336 737 -332
rect 730 -337 737 -336
rect 794 -336 795 -332
rect 799 -336 803 -332
rect 794 -337 803 -336
rect 805 -329 813 -328
rect 805 -333 807 -329
rect 811 -333 813 -329
rect 805 -337 813 -333
rect 815 -331 823 -328
rect 815 -335 817 -331
rect 821 -335 823 -331
rect 815 -337 823 -335
rect 730 -340 735 -337
rect 635 -343 640 -340
rect 591 -344 597 -343
rect 591 -348 592 -344
rect 596 -348 597 -344
rect 591 -349 597 -348
rect 618 -344 624 -343
rect 618 -348 619 -344
rect 623 -348 624 -344
rect 713 -341 719 -340
rect 713 -345 714 -341
rect 718 -345 719 -341
rect 713 -346 719 -345
rect 818 -340 823 -337
rect 825 -340 830 -328
rect 832 -340 840 -328
rect 864 -329 871 -328
rect 866 -332 871 -329
rect 873 -328 878 -323
rect 873 -332 887 -328
rect 878 -336 879 -332
rect 883 -336 887 -332
rect 878 -337 887 -336
rect 889 -329 897 -328
rect 889 -333 891 -329
rect 895 -333 897 -329
rect 889 -337 897 -333
rect 899 -331 907 -328
rect 899 -335 901 -331
rect 905 -335 907 -331
rect 899 -337 907 -335
rect 834 -341 840 -340
rect 834 -345 835 -341
rect 839 -345 840 -341
rect 834 -346 840 -345
rect 902 -340 907 -337
rect 909 -340 914 -328
rect 916 -340 924 -328
rect 934 -329 941 -328
rect 934 -333 935 -329
rect 939 -333 941 -329
rect 934 -334 941 -333
rect 943 -331 951 -328
rect 1692 -307 1704 -305
rect 1692 -311 1695 -307
rect 1699 -310 1704 -307
rect 1699 -311 1701 -310
rect 1692 -313 1701 -311
rect 1692 -317 1701 -315
rect 1692 -321 1693 -317
rect 1697 -321 1701 -317
rect 1692 -323 1701 -321
rect 943 -334 953 -331
rect 945 -340 953 -334
rect 955 -340 960 -331
rect 962 -332 969 -331
rect 962 -336 964 -332
rect 968 -336 969 -332
rect 962 -337 969 -336
rect 962 -340 967 -337
rect 918 -341 924 -340
rect 918 -345 919 -341
rect 923 -345 924 -341
rect 918 -346 924 -345
rect 945 -341 951 -340
rect 945 -345 946 -341
rect 950 -345 951 -341
rect 945 -346 951 -345
rect 618 -349 624 -348
rect 289 -351 295 -350
rect 795 -363 802 -362
rect 468 -366 475 -365
rect 139 -368 146 -367
rect 139 -372 140 -368
rect 144 -372 146 -368
rect 139 -373 146 -372
rect 148 -368 156 -367
rect 148 -372 150 -368
rect 154 -372 156 -368
rect 148 -373 156 -372
rect 158 -368 166 -367
rect 158 -372 160 -368
rect 164 -372 166 -368
rect 158 -373 166 -372
rect 168 -368 175 -367
rect 168 -372 170 -368
rect 174 -372 175 -368
rect 468 -370 469 -366
rect 473 -370 475 -366
rect 468 -371 475 -370
rect 477 -366 485 -365
rect 477 -370 479 -366
rect 483 -370 485 -366
rect 477 -371 485 -370
rect 487 -366 495 -365
rect 487 -370 489 -366
rect 493 -370 495 -366
rect 487 -371 495 -370
rect 497 -366 504 -365
rect 497 -370 499 -366
rect 503 -370 504 -366
rect 795 -367 796 -363
rect 800 -367 802 -363
rect 795 -368 802 -367
rect 804 -363 812 -362
rect 804 -367 806 -363
rect 810 -367 812 -363
rect 804 -368 812 -367
rect 814 -363 822 -362
rect 814 -367 816 -363
rect 820 -367 822 -363
rect 814 -368 822 -367
rect 824 -363 831 -362
rect 824 -367 826 -363
rect 830 -367 831 -363
rect 824 -368 831 -367
rect 497 -371 504 -370
rect 168 -373 175 -372
rect 1692 -329 1701 -325
rect 1692 -333 1696 -329
rect 1700 -333 1701 -329
rect 1692 -334 1701 -333
rect 1687 -339 1696 -334
rect 1687 -343 1696 -341
rect 1687 -347 1688 -343
rect 1692 -346 1696 -343
rect 1692 -347 1693 -346
rect 1687 -348 1693 -347
rect 1410 -372 1417 -371
rect 1410 -376 1411 -372
rect 1415 -376 1417 -372
rect 1410 -377 1417 -376
rect 1412 -381 1417 -377
rect 1419 -380 1429 -371
rect 1419 -381 1422 -380
rect 1421 -384 1422 -381
rect 1426 -384 1429 -380
rect 1421 -385 1429 -384
rect 1431 -372 1438 -371
rect 1431 -376 1433 -372
rect 1437 -376 1438 -372
rect 1431 -379 1438 -376
rect 1692 -373 1710 -372
rect 1692 -377 1705 -373
rect 1709 -377 1710 -373
rect 1692 -378 1710 -377
rect 1431 -383 1433 -379
rect 1437 -383 1438 -379
rect 1692 -380 1704 -378
rect 1431 -385 1438 -383
rect 1051 -406 1062 -403
rect 1064 -406 1081 -403
rect 1726 -382 1732 -381
rect 1692 -387 1704 -382
rect 1692 -391 1704 -389
rect 1692 -395 1695 -391
rect 1699 -394 1704 -391
rect 1699 -395 1701 -394
rect 1692 -397 1701 -395
rect 1163 -402 1173 -401
rect 1123 -407 1134 -404
rect 1136 -407 1153 -404
rect 1163 -406 1165 -402
rect 1169 -406 1173 -402
rect 1163 -407 1173 -406
rect 1175 -407 1194 -401
rect 1196 -402 1204 -401
rect 1196 -406 1199 -402
rect 1203 -406 1204 -402
rect 1196 -407 1204 -406
rect 1217 -402 1227 -401
rect 1217 -406 1219 -402
rect 1223 -406 1227 -402
rect 1217 -407 1227 -406
rect 1229 -407 1248 -401
rect 1250 -402 1258 -401
rect 1250 -406 1253 -402
rect 1257 -406 1258 -402
rect 1250 -407 1258 -406
rect 1273 -402 1283 -401
rect 1273 -406 1275 -402
rect 1279 -406 1283 -402
rect 1273 -407 1283 -406
rect 1285 -407 1304 -401
rect 1306 -402 1314 -401
rect 1306 -406 1309 -402
rect 1313 -406 1314 -402
rect 1306 -407 1314 -406
rect 1327 -402 1337 -401
rect 1327 -406 1329 -402
rect 1333 -406 1337 -402
rect 1327 -407 1337 -406
rect 1339 -407 1358 -401
rect 1360 -402 1368 -401
rect 1360 -406 1363 -402
rect 1367 -406 1368 -402
rect 1360 -407 1368 -406
rect 1692 -401 1701 -399
rect 1692 -405 1693 -401
rect 1697 -405 1701 -401
rect 1692 -407 1701 -405
rect 1692 -413 1701 -409
rect 1127 -429 1138 -426
rect 1140 -429 1157 -426
rect 1167 -427 1177 -426
rect 1167 -431 1169 -427
rect 1173 -431 1177 -427
rect 1167 -432 1177 -431
rect 1179 -432 1198 -426
rect 1200 -427 1208 -426
rect 1200 -431 1203 -427
rect 1207 -431 1208 -427
rect 1200 -432 1208 -431
rect 1221 -427 1231 -426
rect 1221 -431 1223 -427
rect 1227 -431 1231 -427
rect 1221 -432 1231 -431
rect 1233 -432 1252 -426
rect 1254 -427 1262 -426
rect 1254 -431 1257 -427
rect 1261 -431 1262 -427
rect 1254 -432 1262 -431
rect 1277 -427 1287 -426
rect 1277 -431 1279 -427
rect 1283 -431 1287 -427
rect 1277 -432 1287 -431
rect 1289 -432 1308 -426
rect 1310 -427 1318 -426
rect 1310 -431 1313 -427
rect 1317 -431 1318 -427
rect 1310 -432 1318 -431
rect 1331 -427 1341 -426
rect 1331 -431 1333 -427
rect 1337 -431 1341 -427
rect 1331 -432 1341 -431
rect 1343 -432 1362 -426
rect 1364 -427 1372 -426
rect 1423 -424 1431 -423
rect 1423 -427 1424 -424
rect 1364 -431 1367 -427
rect 1371 -431 1372 -427
rect 1414 -431 1419 -427
rect 1364 -432 1372 -431
rect 1412 -432 1419 -431
rect 1412 -436 1413 -432
rect 1417 -436 1419 -432
rect 1412 -437 1419 -436
rect 1421 -428 1424 -427
rect 1428 -428 1431 -424
rect 1421 -437 1431 -428
rect 1433 -425 1440 -423
rect 1692 -417 1696 -413
rect 1700 -417 1701 -413
rect 1692 -418 1701 -417
rect 1687 -423 1696 -418
rect 1726 -386 1727 -382
rect 1731 -386 1732 -382
rect 1726 -388 1732 -386
rect 1726 -392 1732 -390
rect 1726 -396 1727 -392
rect 1731 -396 1732 -392
rect 1726 -398 1732 -396
rect 1726 -402 1732 -400
rect 1726 -406 1727 -402
rect 1731 -406 1732 -402
rect 1726 -408 1732 -406
rect 1726 -412 1732 -410
rect 1726 -416 1727 -412
rect 1731 -416 1732 -412
rect 1726 -417 1732 -416
rect 1433 -429 1435 -425
rect 1439 -429 1440 -425
rect 1433 -432 1440 -429
rect 1687 -427 1696 -425
rect 1687 -431 1688 -427
rect 1692 -430 1696 -427
rect 1692 -431 1693 -430
rect 1723 -430 1729 -429
rect 1723 -431 1724 -430
rect 1687 -432 1693 -431
rect 1433 -436 1435 -432
rect 1439 -436 1440 -432
rect 1716 -434 1724 -431
rect 1728 -434 1729 -430
rect 1716 -436 1729 -434
rect 1433 -437 1440 -436
rect 1716 -440 1729 -438
rect 1716 -443 1720 -440
rect 1719 -444 1720 -443
rect 1724 -444 1729 -440
rect 1719 -446 1729 -444
rect 342 -481 347 -478
rect 340 -482 347 -481
rect 340 -486 341 -482
rect 345 -486 347 -482
rect 340 -487 347 -486
rect 349 -487 360 -478
rect 351 -489 360 -487
rect 362 -489 367 -478
rect 369 -483 374 -478
rect 435 -481 440 -478
rect 433 -482 440 -481
rect 369 -484 376 -483
rect 369 -488 371 -484
rect 375 -488 376 -484
rect 433 -486 434 -482
rect 438 -486 440 -482
rect 433 -487 440 -486
rect 442 -487 453 -478
rect 369 -489 376 -488
rect 351 -494 358 -489
rect 444 -489 453 -487
rect 455 -489 460 -478
rect 462 -483 467 -478
rect 522 -481 527 -478
rect 520 -482 527 -481
rect 462 -484 469 -483
rect 462 -488 464 -484
rect 468 -488 469 -484
rect 520 -486 521 -482
rect 525 -486 527 -482
rect 520 -487 527 -486
rect 529 -487 540 -478
rect 462 -489 469 -488
rect 351 -498 352 -494
rect 356 -498 358 -494
rect 351 -499 358 -498
rect 444 -494 451 -489
rect 531 -489 540 -487
rect 542 -489 547 -478
rect 549 -483 554 -478
rect 1719 -450 1729 -448
rect 1719 -453 1723 -450
rect 1722 -454 1723 -453
rect 1727 -451 1729 -450
rect 1727 -454 1736 -451
rect 1722 -456 1736 -454
rect 1722 -460 1736 -458
rect 1722 -464 1731 -460
rect 1735 -464 1736 -460
rect 1722 -466 1736 -464
rect 1722 -470 1736 -468
rect 1722 -474 1724 -470
rect 1728 -474 1731 -470
rect 1735 -474 1736 -470
rect 1722 -475 1736 -474
rect 549 -484 556 -483
rect 549 -488 551 -484
rect 555 -488 556 -484
rect 549 -489 556 -488
rect 444 -498 445 -494
rect 449 -498 451 -494
rect 444 -499 451 -498
rect 531 -494 538 -489
rect 1695 -476 1701 -475
rect 1695 -480 1696 -476
rect 1700 -477 1701 -476
rect 1700 -480 1704 -477
rect 1695 -482 1704 -480
rect 1723 -480 1729 -479
rect 1723 -481 1724 -480
rect 1716 -484 1724 -481
rect 1728 -481 1729 -480
rect 1728 -484 1736 -481
rect 1695 -489 1704 -484
rect 1716 -486 1736 -484
rect 1695 -493 1704 -491
rect 1716 -493 1736 -488
rect 531 -498 532 -494
rect 536 -498 538 -494
rect 531 -499 538 -498
rect 1692 -494 1710 -493
rect 1692 -498 1705 -494
rect 1709 -498 1710 -494
rect 1692 -499 1710 -498
rect 1716 -497 1736 -495
rect 1692 -501 1698 -499
rect 1716 -501 1717 -497
rect 1721 -501 1736 -497
rect 1716 -502 1736 -501
rect 1692 -505 1698 -503
rect 1692 -509 1693 -505
rect 1697 -509 1698 -505
rect 1716 -504 1730 -502
rect 1716 -508 1730 -506
rect 1692 -510 1698 -509
rect 1716 -511 1724 -508
rect 1723 -512 1724 -511
rect 1728 -512 1730 -508
rect 1723 -513 1730 -512
<< pdiffusion >>
rect 1671 473 1681 474
rect 1671 469 1672 473
rect 1676 469 1681 473
rect 1671 467 1681 469
rect 1671 463 1681 465
rect 1671 459 1676 463
rect 1680 459 1681 463
rect 1671 457 1681 459
rect 1011 433 1042 434
rect 1011 429 1016 433
rect 1020 429 1042 433
rect 1011 428 1042 429
rect 1044 429 1060 434
rect 1605 444 1611 445
rect 1671 453 1681 455
rect 1669 449 1676 453
rect 1680 449 1681 453
rect 1669 447 1681 449
rect 1605 440 1606 444
rect 1610 443 1611 444
rect 1610 440 1617 443
rect 1605 438 1617 440
rect 1669 443 1681 445
rect 1669 440 1676 443
rect 1675 439 1676 440
rect 1680 439 1681 443
rect 1066 429 1079 434
rect 1044 428 1079 429
rect 1099 433 1114 434
rect 1103 429 1114 433
rect 1099 428 1114 429
rect 1116 433 1136 434
rect 1116 429 1132 433
rect 1116 428 1136 429
rect 1143 433 1153 434
rect 1143 429 1145 433
rect 1149 429 1153 433
rect 1143 428 1153 429
rect 1155 433 1174 434
rect 1155 429 1162 433
rect 1166 429 1174 433
rect 1155 428 1174 429
rect 1176 433 1184 434
rect 1176 429 1179 433
rect 1183 429 1184 433
rect 1176 428 1184 429
rect 1197 433 1207 434
rect 1197 429 1199 433
rect 1203 429 1207 433
rect 1197 428 1207 429
rect 1209 433 1228 434
rect 1209 429 1216 433
rect 1220 429 1228 433
rect 1209 428 1228 429
rect 1230 433 1238 434
rect 1230 429 1233 433
rect 1237 429 1238 433
rect 1230 428 1238 429
rect 1253 433 1263 434
rect 1253 429 1255 433
rect 1259 429 1263 433
rect 1253 428 1263 429
rect 1265 433 1284 434
rect 1265 429 1272 433
rect 1276 429 1284 433
rect 1265 428 1284 429
rect 1286 433 1294 434
rect 1286 429 1289 433
rect 1293 429 1294 433
rect 1286 428 1294 429
rect 1307 433 1317 434
rect 1307 429 1309 433
rect 1313 429 1317 433
rect 1307 428 1317 429
rect 1319 433 1338 434
rect 1319 429 1326 433
rect 1330 429 1338 433
rect 1319 428 1338 429
rect 1340 433 1348 434
rect 1340 429 1343 433
rect 1347 429 1348 433
rect 1340 428 1348 429
rect 1605 434 1617 436
rect 1605 430 1606 434
rect 1610 430 1617 434
rect 1605 428 1615 430
rect 1675 438 1681 439
rect 135 403 141 410
rect 114 395 121 403
rect 114 391 115 395
rect 119 391 121 395
rect 114 390 121 391
rect 123 402 131 403
rect 123 398 125 402
rect 129 398 131 402
rect 123 395 131 398
rect 123 391 125 395
rect 129 391 131 395
rect 123 390 131 391
rect 133 397 141 403
rect 133 393 135 397
rect 139 393 141 397
rect 133 392 141 393
rect 143 409 150 410
rect 143 405 145 409
rect 149 405 150 409
rect 143 402 150 405
rect 222 403 228 410
rect 143 398 145 402
rect 149 398 150 402
rect 143 397 150 398
rect 143 392 148 397
rect 201 395 208 403
rect 133 390 139 392
rect 201 391 202 395
rect 206 391 208 395
rect 201 390 208 391
rect 210 402 218 403
rect 210 398 212 402
rect 216 398 218 402
rect 210 395 218 398
rect 210 391 212 395
rect 216 391 218 395
rect 210 390 218 391
rect 220 397 228 403
rect 220 393 222 397
rect 226 393 228 397
rect 220 392 228 393
rect 230 409 237 410
rect 230 405 232 409
rect 236 405 237 409
rect 230 402 237 405
rect 534 411 541 412
rect 315 403 321 410
rect 230 398 232 402
rect 236 398 237 402
rect 230 397 237 398
rect 230 392 235 397
rect 294 395 301 403
rect 220 390 226 392
rect 294 391 295 395
rect 299 391 301 395
rect 294 390 301 391
rect 303 402 311 403
rect 303 398 305 402
rect 309 398 311 402
rect 303 395 311 398
rect 303 391 305 395
rect 309 391 311 395
rect 303 390 311 391
rect 313 397 321 403
rect 313 393 315 397
rect 319 393 321 397
rect 313 392 321 393
rect 323 409 330 410
rect 323 405 325 409
rect 329 405 330 409
rect 323 402 330 405
rect 323 398 325 402
rect 329 398 330 402
rect 534 407 535 411
rect 539 407 541 411
rect 534 404 541 407
rect 534 400 535 404
rect 539 400 541 404
rect 534 399 541 400
rect 323 397 330 398
rect 323 392 328 397
rect 536 394 541 399
rect 543 405 549 412
rect 627 411 634 412
rect 627 407 628 411
rect 632 407 634 411
rect 543 399 551 405
rect 543 395 545 399
rect 549 395 551 399
rect 543 394 551 395
rect 313 390 319 392
rect 545 392 551 394
rect 553 404 561 405
rect 553 400 555 404
rect 559 400 561 404
rect 553 397 561 400
rect 553 393 555 397
rect 559 393 561 397
rect 553 392 561 393
rect 563 397 570 405
rect 627 404 634 407
rect 627 400 628 404
rect 632 400 634 404
rect 627 399 634 400
rect 563 393 565 397
rect 569 393 570 397
rect 629 394 634 399
rect 636 405 642 412
rect 714 411 721 412
rect 714 407 715 411
rect 719 407 721 411
rect 636 399 644 405
rect 636 395 638 399
rect 642 395 644 399
rect 636 394 644 395
rect 563 392 570 393
rect 638 392 644 394
rect 646 404 654 405
rect 646 400 648 404
rect 652 400 654 404
rect 646 397 654 400
rect 646 393 648 397
rect 652 393 654 397
rect 646 392 654 393
rect 656 397 663 405
rect 714 404 721 407
rect 714 400 715 404
rect 719 400 721 404
rect 714 399 721 400
rect 656 393 658 397
rect 662 393 663 397
rect 716 394 721 399
rect 723 405 729 412
rect 1605 424 1615 426
rect 1605 420 1606 424
rect 1610 420 1615 424
rect 1659 427 1665 428
rect 1659 426 1660 427
rect 1605 418 1615 420
rect 723 399 731 405
rect 723 395 725 399
rect 729 395 731 399
rect 723 394 731 395
rect 656 392 663 393
rect 725 392 731 394
rect 733 404 741 405
rect 733 400 735 404
rect 739 400 741 404
rect 733 397 741 400
rect 733 393 735 397
rect 739 393 741 397
rect 733 392 741 393
rect 743 397 750 405
rect 743 393 745 397
rect 749 393 750 397
rect 743 392 750 393
rect 1605 414 1615 416
rect 1605 410 1610 414
rect 1614 410 1615 414
rect 1653 423 1660 426
rect 1664 426 1665 427
rect 1664 423 1680 426
rect 1653 421 1680 423
rect 1653 417 1680 419
rect 1653 414 1668 417
rect 1662 413 1668 414
rect 1672 413 1680 417
rect 1662 411 1680 413
rect 1605 409 1615 410
rect 1662 407 1680 409
rect 1662 403 1675 407
rect 1679 403 1680 407
rect 1662 401 1680 403
rect 1662 397 1680 399
rect 1653 391 1680 397
rect 1653 387 1654 391
rect 1658 387 1661 391
rect 1665 387 1680 391
rect 1653 385 1680 387
rect 1653 381 1680 383
rect 1653 378 1675 381
rect 1674 377 1675 378
rect 1679 377 1680 381
rect 1674 376 1680 377
rect 38 342 43 348
rect 36 341 43 342
rect 36 337 37 341
rect 41 337 43 341
rect 36 336 43 337
rect 45 346 51 348
rect 45 341 53 346
rect 45 337 47 341
rect 51 337 53 341
rect 45 336 53 337
rect 55 341 63 346
rect 55 337 57 341
rect 61 337 63 341
rect 55 336 63 337
rect 65 345 72 346
rect 65 341 67 345
rect 71 341 72 345
rect 124 343 129 364
rect 65 336 72 341
rect 122 342 129 343
rect 122 338 123 342
rect 127 338 129 342
rect 122 337 129 338
rect 131 363 143 364
rect 131 359 133 363
rect 137 359 143 363
rect 131 356 143 359
rect 131 352 133 356
rect 137 355 143 356
rect 160 355 165 364
rect 137 352 145 355
rect 131 337 145 352
rect 147 342 155 355
rect 147 338 149 342
rect 153 338 155 342
rect 147 337 155 338
rect 157 349 165 355
rect 157 345 159 349
rect 163 345 165 349
rect 157 337 165 345
rect 167 358 172 364
rect 167 357 174 358
rect 167 353 169 357
rect 173 353 174 357
rect 167 352 174 353
rect 167 337 172 352
rect 208 343 213 364
rect 206 342 213 343
rect 206 338 207 342
rect 211 338 213 342
rect 206 337 213 338
rect 215 363 227 364
rect 215 359 217 363
rect 221 359 227 363
rect 215 356 227 359
rect 215 352 217 356
rect 221 355 227 356
rect 244 355 249 364
rect 221 352 229 355
rect 215 337 229 352
rect 231 342 239 355
rect 231 338 233 342
rect 237 338 239 342
rect 231 337 239 338
rect 241 349 249 355
rect 241 345 243 349
rect 247 345 249 349
rect 241 337 249 345
rect 251 358 256 364
rect 251 357 258 358
rect 251 353 253 357
rect 257 353 258 357
rect 251 352 258 353
rect 251 337 256 352
rect 270 342 275 348
rect 268 341 275 342
rect 268 337 269 341
rect 273 337 275 341
rect 268 336 275 337
rect 277 346 283 348
rect 277 341 285 346
rect 277 337 279 341
rect 283 337 285 341
rect 277 336 285 337
rect 287 341 295 346
rect 287 337 289 341
rect 293 337 295 341
rect 287 336 295 337
rect 297 345 304 346
rect 297 341 299 345
rect 303 341 304 345
rect 367 344 372 350
rect 297 336 304 341
rect 365 343 372 344
rect 365 339 366 343
rect 370 339 372 343
rect 365 338 372 339
rect 374 348 380 350
rect 374 343 382 348
rect 374 339 376 343
rect 380 339 382 343
rect 374 338 382 339
rect 384 343 392 348
rect 384 339 386 343
rect 390 339 392 343
rect 384 338 392 339
rect 394 347 401 348
rect 394 343 396 347
rect 400 343 401 347
rect 453 345 458 366
rect 394 338 401 343
rect 451 344 458 345
rect 451 340 452 344
rect 456 340 458 344
rect 451 339 458 340
rect 460 365 472 366
rect 460 361 462 365
rect 466 361 472 365
rect 460 358 472 361
rect 460 354 462 358
rect 466 357 472 358
rect 489 357 494 366
rect 466 354 474 357
rect 460 339 474 354
rect 476 344 484 357
rect 476 340 478 344
rect 482 340 484 344
rect 476 339 484 340
rect 486 351 494 357
rect 486 347 488 351
rect 492 347 494 351
rect 486 339 494 347
rect 496 360 501 366
rect 496 359 503 360
rect 496 355 498 359
rect 502 355 503 359
rect 496 354 503 355
rect 496 339 501 354
rect 537 345 542 366
rect 535 344 542 345
rect 535 340 536 344
rect 540 340 542 344
rect 535 339 542 340
rect 544 365 556 366
rect 544 361 546 365
rect 550 361 556 365
rect 544 358 556 361
rect 544 354 546 358
rect 550 357 556 358
rect 573 357 578 366
rect 550 354 558 357
rect 544 339 558 354
rect 560 344 568 357
rect 560 340 562 344
rect 566 340 568 344
rect 560 339 568 340
rect 570 351 578 357
rect 570 347 572 351
rect 576 347 578 351
rect 570 339 578 347
rect 580 360 585 366
rect 580 359 587 360
rect 580 355 582 359
rect 586 355 587 359
rect 580 354 587 355
rect 580 339 585 354
rect 599 344 604 350
rect 597 343 604 344
rect 597 339 598 343
rect 602 339 604 343
rect 597 338 604 339
rect 606 348 612 350
rect 606 343 614 348
rect 606 339 608 343
rect 612 339 614 343
rect 606 338 614 339
rect 616 343 624 348
rect 616 339 618 343
rect 622 339 624 343
rect 616 338 624 339
rect 626 347 633 348
rect 694 347 699 353
rect 626 343 628 347
rect 632 343 633 347
rect 626 338 633 343
rect 692 346 699 347
rect 692 342 693 346
rect 697 342 699 346
rect 692 341 699 342
rect 701 351 707 353
rect 701 346 709 351
rect 701 342 703 346
rect 707 342 709 346
rect 701 341 709 342
rect 711 346 719 351
rect 711 342 713 346
rect 717 342 719 346
rect 711 341 719 342
rect 721 350 728 351
rect 721 346 723 350
rect 727 346 728 350
rect 780 348 785 369
rect 721 341 728 346
rect 778 347 785 348
rect 778 343 779 347
rect 783 343 785 347
rect 778 342 785 343
rect 787 368 799 369
rect 787 364 789 368
rect 793 364 799 368
rect 787 361 799 364
rect 787 357 789 361
rect 793 360 799 361
rect 816 360 821 369
rect 793 357 801 360
rect 787 342 801 357
rect 803 347 811 360
rect 803 343 805 347
rect 809 343 811 347
rect 803 342 811 343
rect 813 354 821 360
rect 813 350 815 354
rect 819 350 821 354
rect 813 342 821 350
rect 823 363 828 369
rect 823 362 830 363
rect 823 358 825 362
rect 829 358 830 362
rect 823 357 830 358
rect 823 342 828 357
rect 864 348 869 369
rect 862 347 869 348
rect 862 343 863 347
rect 867 343 869 347
rect 862 342 869 343
rect 871 368 883 369
rect 871 364 873 368
rect 877 364 883 368
rect 871 361 883 364
rect 871 357 873 361
rect 877 360 883 361
rect 900 360 905 369
rect 877 357 885 360
rect 871 342 885 357
rect 887 347 895 360
rect 887 343 889 347
rect 893 343 895 347
rect 887 342 895 343
rect 897 354 905 360
rect 897 350 899 354
rect 903 350 905 354
rect 897 342 905 350
rect 907 363 912 369
rect 907 362 914 363
rect 907 358 909 362
rect 913 358 914 362
rect 907 357 914 358
rect 907 342 912 357
rect 926 347 931 353
rect 924 346 931 347
rect 924 342 925 346
rect 929 342 931 346
rect 924 341 931 342
rect 933 351 939 353
rect 933 346 941 351
rect 933 342 935 346
rect 939 342 941 346
rect 933 341 941 342
rect 943 346 951 351
rect 943 342 945 346
rect 949 342 951 346
rect 943 341 951 342
rect 953 350 960 351
rect 953 346 955 350
rect 959 346 960 350
rect 1510 351 1516 352
rect 1510 350 1511 351
rect 953 341 960 346
rect 1503 347 1511 350
rect 1515 350 1516 351
rect 1515 347 1521 350
rect 1503 345 1521 347
rect 1503 338 1521 343
rect 1103 334 1118 335
rect 1107 330 1118 334
rect 1103 329 1118 330
rect 1120 334 1140 335
rect 1120 330 1136 334
rect 1120 329 1140 330
rect 1147 334 1157 335
rect 1147 330 1149 334
rect 1153 330 1157 334
rect 1147 329 1157 330
rect 1159 334 1178 335
rect 1159 330 1166 334
rect 1170 330 1178 334
rect 1159 329 1178 330
rect 1180 334 1188 335
rect 1180 330 1183 334
rect 1187 330 1188 334
rect 1180 329 1188 330
rect 1201 334 1211 335
rect 1201 330 1203 334
rect 1207 330 1211 334
rect 1201 329 1211 330
rect 1213 334 1232 335
rect 1213 330 1220 334
rect 1224 330 1232 334
rect 1213 329 1232 330
rect 1234 334 1242 335
rect 1234 330 1237 334
rect 1241 330 1242 334
rect 1234 329 1242 330
rect 1257 334 1267 335
rect 1257 330 1259 334
rect 1263 330 1267 334
rect 1257 329 1267 330
rect 1269 334 1288 335
rect 1269 330 1276 334
rect 1280 330 1288 334
rect 1269 329 1288 330
rect 1290 334 1298 335
rect 1290 330 1293 334
rect 1297 330 1298 334
rect 1290 329 1298 330
rect 1311 334 1321 335
rect 1311 330 1313 334
rect 1317 330 1321 334
rect 1311 329 1321 330
rect 1323 334 1342 335
rect 1323 330 1330 334
rect 1334 330 1342 334
rect 1323 329 1342 330
rect 1344 334 1352 335
rect 1344 330 1347 334
rect 1351 330 1352 334
rect 1344 329 1352 330
rect 1503 333 1521 336
rect 1503 329 1504 333
rect 1508 329 1524 333
rect 1503 327 1524 329
rect 1512 325 1524 327
rect 1512 321 1524 323
rect 1512 317 1513 321
rect 1517 318 1524 321
rect 1517 317 1518 318
rect 1512 316 1518 317
rect 1606 358 1612 359
rect 1606 354 1607 358
rect 1611 357 1612 358
rect 1611 354 1633 357
rect 1606 352 1633 354
rect 1606 348 1633 350
rect 1606 344 1621 348
rect 1625 344 1628 348
rect 1632 344 1633 348
rect 1606 338 1633 344
rect 1659 343 1665 344
rect 1659 342 1660 343
rect 1653 339 1660 342
rect 1664 342 1665 343
rect 1664 339 1680 342
rect 1606 336 1624 338
rect 1653 337 1680 339
rect 1606 332 1624 334
rect 1653 333 1680 335
rect 1606 328 1607 332
rect 1611 328 1624 332
rect 1606 326 1624 328
rect 1653 330 1668 333
rect 1662 329 1668 330
rect 1672 329 1680 333
rect 1662 327 1680 329
rect 1606 322 1624 324
rect 1606 318 1614 322
rect 1618 321 1624 322
rect 1618 318 1633 321
rect 1662 323 1680 325
rect 1662 319 1675 323
rect 1679 319 1680 323
rect 1606 316 1633 318
rect 1662 317 1680 319
rect 1606 312 1633 314
rect 1662 313 1680 315
rect 1606 309 1622 312
rect 1387 306 1393 307
rect 1387 302 1388 306
rect 1392 304 1393 306
rect 1621 308 1622 309
rect 1626 309 1633 312
rect 1626 308 1627 309
rect 1621 307 1627 308
rect 1653 307 1680 313
rect 1392 302 1395 304
rect 1011 288 1042 289
rect 1011 284 1016 288
rect 1020 284 1042 288
rect 148 252 156 255
rect 131 247 136 252
rect 129 246 136 247
rect 129 242 130 246
rect 134 242 136 246
rect 129 241 136 242
rect 131 234 136 241
rect 138 234 143 252
rect 145 243 156 252
rect 158 249 163 255
rect 1011 283 1042 284
rect 1044 284 1060 289
rect 1387 293 1395 302
rect 1378 289 1383 293
rect 1066 284 1079 289
rect 1044 283 1079 284
rect 1099 288 1114 289
rect 1103 284 1114 288
rect 1099 283 1114 284
rect 1116 288 1136 289
rect 1116 284 1132 288
rect 1116 283 1136 284
rect 1143 288 1153 289
rect 1143 284 1145 288
rect 1149 284 1153 288
rect 1143 283 1153 284
rect 1155 288 1174 289
rect 1155 284 1162 288
rect 1166 284 1174 288
rect 1155 283 1174 284
rect 1176 288 1184 289
rect 1176 284 1179 288
rect 1183 284 1184 288
rect 1176 283 1184 284
rect 1197 288 1207 289
rect 1197 284 1199 288
rect 1203 284 1207 288
rect 1197 283 1207 284
rect 1209 288 1228 289
rect 1209 284 1216 288
rect 1220 284 1228 288
rect 1209 283 1228 284
rect 1230 288 1238 289
rect 1230 284 1233 288
rect 1237 284 1238 288
rect 1230 283 1238 284
rect 1253 288 1263 289
rect 1253 284 1255 288
rect 1259 284 1263 288
rect 1253 283 1263 284
rect 1265 288 1284 289
rect 1265 284 1272 288
rect 1276 284 1284 288
rect 1265 283 1284 284
rect 1286 288 1294 289
rect 1286 284 1289 288
rect 1293 284 1294 288
rect 1286 283 1294 284
rect 1307 288 1317 289
rect 1307 284 1309 288
rect 1313 284 1317 288
rect 1307 283 1317 284
rect 1319 288 1338 289
rect 1319 284 1326 288
rect 1330 284 1338 288
rect 1319 283 1338 284
rect 1340 288 1348 289
rect 1340 284 1343 288
rect 1347 284 1348 288
rect 1340 283 1348 284
rect 1376 288 1383 289
rect 1376 284 1377 288
rect 1381 284 1383 288
rect 1376 283 1383 284
rect 1378 276 1383 283
rect 1385 276 1395 293
rect 1397 297 1402 304
rect 1653 303 1654 307
rect 1658 303 1661 307
rect 1665 303 1680 307
rect 1653 301 1680 303
rect 1653 297 1680 299
rect 1397 296 1404 297
rect 1397 292 1399 296
rect 1403 292 1404 296
rect 1653 294 1675 297
rect 1674 293 1675 294
rect 1679 293 1680 297
rect 1674 292 1680 293
rect 1768 334 1774 335
rect 1768 333 1769 334
rect 1762 330 1769 333
rect 1773 330 1774 334
rect 1762 328 1774 330
rect 1762 324 1774 326
rect 1762 322 1783 324
rect 1762 318 1778 322
rect 1782 318 1783 322
rect 1765 315 1783 318
rect 1765 308 1783 313
rect 1765 304 1783 306
rect 1765 301 1771 304
rect 1770 300 1771 301
rect 1775 301 1783 304
rect 1775 300 1776 301
rect 1770 299 1776 300
rect 1397 289 1404 292
rect 1397 285 1399 289
rect 1403 285 1404 289
rect 1397 284 1404 285
rect 1397 276 1402 284
rect 804 257 812 260
rect 477 254 485 257
rect 460 249 465 254
rect 158 248 165 249
rect 158 244 160 248
rect 164 244 165 248
rect 158 243 165 244
rect 458 248 465 249
rect 458 244 459 248
rect 463 244 465 248
rect 458 243 465 244
rect 145 239 154 243
rect 145 235 148 239
rect 152 235 154 239
rect 145 234 154 235
rect 460 236 465 243
rect 467 236 472 254
rect 474 245 485 254
rect 487 251 492 257
rect 787 252 792 257
rect 785 251 792 252
rect 487 250 494 251
rect 487 246 489 250
rect 493 246 494 250
rect 785 247 786 251
rect 790 247 792 251
rect 785 246 792 247
rect 487 245 494 246
rect 474 241 483 245
rect 474 237 477 241
rect 481 237 483 241
rect 787 239 792 246
rect 794 239 799 257
rect 801 248 812 257
rect 814 254 819 260
rect 814 253 821 254
rect 814 249 816 253
rect 820 249 821 253
rect 814 248 821 249
rect 801 244 810 248
rect 1606 274 1612 275
rect 1606 270 1607 274
rect 1611 273 1612 274
rect 1611 270 1633 273
rect 1606 268 1633 270
rect 1606 264 1633 266
rect 1606 260 1621 264
rect 1625 260 1628 264
rect 1632 260 1633 264
rect 1606 254 1633 260
rect 1606 252 1624 254
rect 801 240 804 244
rect 808 240 810 244
rect 1606 248 1624 250
rect 801 239 810 240
rect 474 236 483 237
rect 1606 244 1607 248
rect 1611 244 1624 248
rect 1606 242 1624 244
rect 1671 241 1681 242
rect 1606 238 1624 240
rect 37 196 42 202
rect 35 195 42 196
rect 35 191 36 195
rect 40 191 42 195
rect 35 190 42 191
rect 44 200 50 202
rect 44 195 52 200
rect 44 191 46 195
rect 50 191 52 195
rect 44 190 52 191
rect 54 195 62 200
rect 54 191 56 195
rect 60 191 62 195
rect 54 190 62 191
rect 64 199 71 200
rect 64 195 66 199
rect 70 195 71 199
rect 123 197 128 218
rect 64 190 71 195
rect 121 196 128 197
rect 121 192 122 196
rect 126 192 128 196
rect 121 191 128 192
rect 130 217 142 218
rect 130 213 132 217
rect 136 213 142 217
rect 130 210 142 213
rect 130 206 132 210
rect 136 209 142 210
rect 159 209 164 218
rect 136 206 144 209
rect 130 191 144 206
rect 146 196 154 209
rect 146 192 148 196
rect 152 192 154 196
rect 146 191 154 192
rect 156 203 164 209
rect 156 199 158 203
rect 162 199 164 203
rect 156 191 164 199
rect 166 212 171 218
rect 166 211 173 212
rect 166 207 168 211
rect 172 207 173 211
rect 166 206 173 207
rect 166 191 171 206
rect 207 197 212 218
rect 205 196 212 197
rect 205 192 206 196
rect 210 192 212 196
rect 205 191 212 192
rect 214 217 226 218
rect 214 213 216 217
rect 220 213 226 217
rect 214 210 226 213
rect 214 206 216 210
rect 220 209 226 210
rect 243 209 248 218
rect 220 206 228 209
rect 214 191 228 206
rect 230 196 238 209
rect 230 192 232 196
rect 236 192 238 196
rect 230 191 238 192
rect 240 203 248 209
rect 240 199 242 203
rect 246 199 248 203
rect 240 191 248 199
rect 250 212 255 218
rect 250 211 257 212
rect 250 207 252 211
rect 256 207 257 211
rect 250 206 257 207
rect 250 191 255 206
rect 269 196 274 202
rect 267 195 274 196
rect 267 191 268 195
rect 272 191 274 195
rect 267 190 274 191
rect 276 200 282 202
rect 276 195 284 200
rect 276 191 278 195
rect 282 191 284 195
rect 276 190 284 191
rect 286 195 294 200
rect 286 191 288 195
rect 292 191 294 195
rect 286 190 294 191
rect 296 199 303 200
rect 296 195 298 199
rect 302 195 303 199
rect 366 198 371 204
rect 296 190 303 195
rect 364 197 371 198
rect 364 193 365 197
rect 369 193 371 197
rect 364 192 371 193
rect 373 202 379 204
rect 373 197 381 202
rect 373 193 375 197
rect 379 193 381 197
rect 373 192 381 193
rect 383 197 391 202
rect 383 193 385 197
rect 389 193 391 197
rect 383 192 391 193
rect 393 201 400 202
rect 393 197 395 201
rect 399 197 400 201
rect 452 199 457 220
rect 393 192 400 197
rect 450 198 457 199
rect 450 194 451 198
rect 455 194 457 198
rect 450 193 457 194
rect 459 219 471 220
rect 459 215 461 219
rect 465 215 471 219
rect 459 212 471 215
rect 459 208 461 212
rect 465 211 471 212
rect 488 211 493 220
rect 465 208 473 211
rect 459 193 473 208
rect 475 198 483 211
rect 475 194 477 198
rect 481 194 483 198
rect 475 193 483 194
rect 485 205 493 211
rect 485 201 487 205
rect 491 201 493 205
rect 485 193 493 201
rect 495 214 500 220
rect 495 213 502 214
rect 495 209 497 213
rect 501 209 502 213
rect 495 208 502 209
rect 495 193 500 208
rect 536 199 541 220
rect 534 198 541 199
rect 534 194 535 198
rect 539 194 541 198
rect 534 193 541 194
rect 543 219 555 220
rect 543 215 545 219
rect 549 215 555 219
rect 543 212 555 215
rect 543 208 545 212
rect 549 211 555 212
rect 572 211 577 220
rect 549 208 557 211
rect 543 193 557 208
rect 559 198 567 211
rect 559 194 561 198
rect 565 194 567 198
rect 559 193 567 194
rect 569 205 577 211
rect 569 201 571 205
rect 575 201 577 205
rect 569 193 577 201
rect 579 214 584 220
rect 579 213 586 214
rect 579 209 581 213
rect 585 209 586 213
rect 579 208 586 209
rect 579 193 584 208
rect 598 198 603 204
rect 596 197 603 198
rect 596 193 597 197
rect 601 193 603 197
rect 596 192 603 193
rect 605 202 611 204
rect 605 197 613 202
rect 605 193 607 197
rect 611 193 613 197
rect 605 192 613 193
rect 615 197 623 202
rect 615 193 617 197
rect 621 193 623 197
rect 615 192 623 193
rect 625 201 632 202
rect 693 201 698 207
rect 625 197 627 201
rect 631 197 632 201
rect 625 192 632 197
rect 691 200 698 201
rect 691 196 692 200
rect 696 196 698 200
rect 691 195 698 196
rect 700 205 706 207
rect 700 200 708 205
rect 700 196 702 200
rect 706 196 708 200
rect 700 195 708 196
rect 710 200 718 205
rect 710 196 712 200
rect 716 196 718 200
rect 710 195 718 196
rect 720 204 727 205
rect 720 200 722 204
rect 726 200 727 204
rect 779 202 784 223
rect 720 195 727 200
rect 777 201 784 202
rect 777 197 778 201
rect 782 197 784 201
rect 777 196 784 197
rect 786 222 798 223
rect 786 218 788 222
rect 792 218 798 222
rect 786 215 798 218
rect 786 211 788 215
rect 792 214 798 215
rect 815 214 820 223
rect 792 211 800 214
rect 786 196 800 211
rect 802 201 810 214
rect 802 197 804 201
rect 808 197 810 201
rect 802 196 810 197
rect 812 208 820 214
rect 812 204 814 208
rect 818 204 820 208
rect 812 196 820 204
rect 822 217 827 223
rect 822 216 829 217
rect 822 212 824 216
rect 828 212 829 216
rect 822 211 829 212
rect 822 196 827 211
rect 863 202 868 223
rect 861 201 868 202
rect 861 197 862 201
rect 866 197 868 201
rect 861 196 868 197
rect 870 222 882 223
rect 870 218 872 222
rect 876 218 882 222
rect 870 215 882 218
rect 870 211 872 215
rect 876 214 882 215
rect 899 214 904 223
rect 876 211 884 214
rect 870 196 884 211
rect 886 201 894 214
rect 886 197 888 201
rect 892 197 894 201
rect 886 196 894 197
rect 896 208 904 214
rect 896 204 898 208
rect 902 204 904 208
rect 896 196 904 204
rect 906 217 911 223
rect 906 216 913 217
rect 906 212 908 216
rect 912 212 913 216
rect 906 211 913 212
rect 906 196 911 211
rect 925 201 930 207
rect 923 200 930 201
rect 923 196 924 200
rect 928 196 930 200
rect 923 195 930 196
rect 932 205 938 207
rect 1606 234 1614 238
rect 1618 237 1624 238
rect 1618 234 1633 237
rect 1606 232 1633 234
rect 1606 228 1633 230
rect 1606 225 1622 228
rect 1621 224 1622 225
rect 1626 225 1633 228
rect 1671 237 1672 241
rect 1676 237 1681 241
rect 1671 235 1681 237
rect 1671 231 1681 233
rect 1626 224 1627 225
rect 1621 223 1627 224
rect 1671 227 1676 231
rect 1680 227 1681 231
rect 1671 225 1681 227
rect 1605 212 1611 213
rect 1671 221 1681 223
rect 1669 217 1676 221
rect 1680 217 1681 221
rect 1669 215 1681 217
rect 1605 208 1606 212
rect 1610 211 1611 212
rect 1610 208 1617 211
rect 1605 206 1617 208
rect 1669 211 1681 213
rect 1669 208 1676 211
rect 1675 207 1676 208
rect 1680 207 1681 211
rect 932 200 940 205
rect 932 196 934 200
rect 938 196 940 200
rect 932 195 940 196
rect 942 200 950 205
rect 942 196 944 200
rect 948 196 950 200
rect 942 195 950 196
rect 952 204 959 205
rect 952 200 954 204
rect 958 200 959 204
rect 952 195 959 200
rect 1379 196 1384 203
rect 1377 195 1384 196
rect 1377 191 1378 195
rect 1382 191 1384 195
rect 1377 190 1384 191
rect 1103 189 1118 190
rect 1107 185 1118 189
rect 1103 184 1118 185
rect 1120 189 1140 190
rect 1120 185 1136 189
rect 1120 184 1140 185
rect 1147 189 1157 190
rect 1147 185 1149 189
rect 1153 185 1157 189
rect 1147 184 1157 185
rect 1159 189 1178 190
rect 1159 185 1166 189
rect 1170 185 1178 189
rect 1159 184 1178 185
rect 1180 189 1188 190
rect 1180 185 1183 189
rect 1187 185 1188 189
rect 1180 184 1188 185
rect 1201 189 1211 190
rect 1201 185 1203 189
rect 1207 185 1211 189
rect 1201 184 1211 185
rect 1213 189 1232 190
rect 1213 185 1220 189
rect 1224 185 1232 189
rect 1213 184 1232 185
rect 1234 189 1242 190
rect 1234 185 1237 189
rect 1241 185 1242 189
rect 1234 184 1242 185
rect 1257 189 1267 190
rect 1257 185 1259 189
rect 1263 185 1267 189
rect 1257 184 1267 185
rect 1269 189 1288 190
rect 1269 185 1276 189
rect 1280 185 1288 189
rect 1269 184 1288 185
rect 1290 189 1298 190
rect 1290 185 1293 189
rect 1297 185 1298 189
rect 1290 184 1298 185
rect 1311 189 1321 190
rect 1311 185 1313 189
rect 1317 185 1321 189
rect 1311 184 1321 185
rect 1323 189 1342 190
rect 1323 185 1330 189
rect 1334 185 1342 189
rect 1323 184 1342 185
rect 1344 189 1352 190
rect 1344 185 1347 189
rect 1351 185 1352 189
rect 1379 186 1384 190
rect 1386 186 1396 203
rect 1344 184 1352 185
rect 1388 177 1396 186
rect 1388 173 1389 177
rect 1393 175 1396 177
rect 1398 195 1403 203
rect 1605 202 1617 204
rect 1605 198 1606 202
rect 1610 198 1617 202
rect 1605 196 1615 198
rect 1675 206 1681 207
rect 1398 194 1405 195
rect 1398 190 1400 194
rect 1404 190 1405 194
rect 1605 192 1615 194
rect 1398 187 1405 190
rect 1605 188 1606 192
rect 1610 188 1615 192
rect 1398 183 1400 187
rect 1404 183 1405 187
rect 1605 186 1615 188
rect 1398 182 1405 183
rect 1398 175 1403 182
rect 1605 182 1615 184
rect 1605 178 1610 182
rect 1614 178 1615 182
rect 1605 177 1615 178
rect 1393 173 1394 175
rect 1388 172 1394 173
rect 1387 166 1393 167
rect 1387 162 1388 166
rect 1392 164 1393 166
rect 1392 162 1395 164
rect 1387 153 1395 162
rect 1010 146 1041 147
rect 1010 142 1015 146
rect 1019 142 1041 146
rect 1010 141 1041 142
rect 1043 142 1059 147
rect 1378 149 1383 153
rect 1376 148 1383 149
rect 1065 142 1078 147
rect 1043 141 1078 142
rect 1098 146 1113 147
rect 1102 142 1113 146
rect 1098 141 1113 142
rect 1115 146 1135 147
rect 1115 142 1131 146
rect 1115 141 1135 142
rect 1142 146 1152 147
rect 1142 142 1144 146
rect 1148 142 1152 146
rect 1142 141 1152 142
rect 1154 146 1173 147
rect 1154 142 1161 146
rect 1165 142 1173 146
rect 1154 141 1173 142
rect 1175 146 1183 147
rect 1175 142 1178 146
rect 1182 142 1183 146
rect 1175 141 1183 142
rect 1196 146 1206 147
rect 1196 142 1198 146
rect 1202 142 1206 146
rect 1196 141 1206 142
rect 1208 146 1227 147
rect 1208 142 1215 146
rect 1219 142 1227 146
rect 1208 141 1227 142
rect 1229 146 1237 147
rect 1229 142 1232 146
rect 1236 142 1237 146
rect 1229 141 1237 142
rect 1252 146 1262 147
rect 1252 142 1254 146
rect 1258 142 1262 146
rect 1252 141 1262 142
rect 1264 146 1283 147
rect 1264 142 1271 146
rect 1275 142 1283 146
rect 1264 141 1283 142
rect 1285 146 1293 147
rect 1285 142 1288 146
rect 1292 142 1293 146
rect 1285 141 1293 142
rect 1306 146 1316 147
rect 1306 142 1308 146
rect 1312 142 1316 146
rect 1306 141 1316 142
rect 1318 146 1337 147
rect 1318 142 1325 146
rect 1329 142 1337 146
rect 1318 141 1337 142
rect 1339 146 1347 147
rect 1339 142 1342 146
rect 1346 142 1347 146
rect 1376 144 1377 148
rect 1381 144 1383 148
rect 1376 143 1383 144
rect 1339 141 1347 142
rect 147 106 155 109
rect 130 101 135 106
rect 128 100 135 101
rect 128 96 129 100
rect 133 96 135 100
rect 128 95 135 96
rect 130 88 135 95
rect 137 88 142 106
rect 144 97 155 106
rect 157 103 162 109
rect 1378 136 1383 143
rect 1385 136 1395 153
rect 1397 157 1402 164
rect 1397 156 1404 157
rect 1397 152 1399 156
rect 1403 152 1404 156
rect 1397 149 1404 152
rect 1397 145 1399 149
rect 1403 145 1404 149
rect 1397 144 1404 145
rect 1397 136 1402 144
rect 803 111 811 114
rect 476 108 484 111
rect 459 103 464 108
rect 157 102 164 103
rect 157 98 159 102
rect 163 98 164 102
rect 157 97 164 98
rect 457 102 464 103
rect 457 98 458 102
rect 462 98 464 102
rect 457 97 464 98
rect 144 93 153 97
rect 144 89 147 93
rect 151 89 153 93
rect 144 88 153 89
rect 459 90 464 97
rect 466 90 471 108
rect 473 99 484 108
rect 486 105 491 111
rect 786 106 791 111
rect 784 105 791 106
rect 486 104 493 105
rect 486 100 488 104
rect 492 100 493 104
rect 784 101 785 105
rect 789 101 791 105
rect 784 100 791 101
rect 486 99 493 100
rect 473 95 482 99
rect 473 91 476 95
rect 480 91 482 95
rect 786 93 791 100
rect 793 93 798 111
rect 800 102 811 111
rect 813 108 818 114
rect 813 107 820 108
rect 813 103 815 107
rect 819 103 820 107
rect 813 102 820 103
rect 1673 113 1683 114
rect 800 98 809 102
rect 1673 109 1674 113
rect 1678 109 1683 113
rect 1673 107 1683 109
rect 1673 103 1683 105
rect 800 94 803 98
rect 807 94 809 98
rect 800 93 809 94
rect 473 90 482 91
rect 1673 99 1678 103
rect 1682 99 1683 103
rect 1673 97 1683 99
rect 340 61 346 63
rect 331 56 336 61
rect 329 55 336 56
rect 329 51 330 55
rect 334 51 336 55
rect 329 48 336 51
rect 329 44 330 48
rect 334 44 336 48
rect 329 43 336 44
rect 338 60 346 61
rect 338 56 340 60
rect 344 56 346 60
rect 338 50 346 56
rect 348 62 356 63
rect 348 58 350 62
rect 354 58 356 62
rect 348 55 356 58
rect 348 51 350 55
rect 354 51 356 55
rect 348 50 356 51
rect 358 62 365 63
rect 358 58 360 62
rect 364 58 365 62
rect 433 61 439 63
rect 358 50 365 58
rect 424 56 429 61
rect 422 55 429 56
rect 422 51 423 55
rect 427 51 429 55
rect 338 43 344 50
rect 422 48 429 51
rect 422 44 423 48
rect 427 44 429 48
rect 422 43 429 44
rect 431 60 439 61
rect 431 56 433 60
rect 437 56 439 60
rect 431 50 439 56
rect 441 62 449 63
rect 441 58 443 62
rect 447 58 449 62
rect 441 55 449 58
rect 441 51 443 55
rect 447 51 449 55
rect 441 50 449 51
rect 451 62 458 63
rect 451 58 453 62
rect 457 58 458 62
rect 1607 84 1613 85
rect 1673 93 1683 95
rect 1671 89 1678 93
rect 1682 89 1683 93
rect 1671 87 1683 89
rect 1607 80 1608 84
rect 1612 83 1613 84
rect 1612 80 1619 83
rect 1607 78 1619 80
rect 1671 83 1683 85
rect 1671 80 1678 83
rect 1677 79 1678 80
rect 1682 79 1683 83
rect 1607 74 1619 76
rect 1607 70 1608 74
rect 1612 70 1619 74
rect 1607 68 1617 70
rect 1677 78 1683 79
rect 1607 64 1617 66
rect 520 61 526 63
rect 451 50 458 58
rect 511 56 516 61
rect 509 55 516 56
rect 509 51 510 55
rect 514 51 516 55
rect 431 43 437 50
rect 509 48 516 51
rect 509 44 510 48
rect 514 44 516 48
rect 509 43 516 44
rect 518 60 526 61
rect 518 56 520 60
rect 524 56 526 60
rect 518 50 526 56
rect 528 62 536 63
rect 528 58 530 62
rect 534 58 536 62
rect 528 55 536 58
rect 528 51 530 55
rect 534 51 536 55
rect 528 50 536 51
rect 538 62 545 63
rect 538 58 540 62
rect 544 58 545 62
rect 538 50 545 58
rect 518 43 524 50
rect 1607 60 1608 64
rect 1612 60 1617 64
rect 1661 67 1667 68
rect 1661 66 1662 67
rect 1607 58 1617 60
rect 1607 54 1617 56
rect 1607 50 1612 54
rect 1616 50 1617 54
rect 1655 63 1662 66
rect 1666 66 1667 67
rect 1666 63 1682 66
rect 1655 61 1682 63
rect 1655 57 1682 59
rect 1655 54 1670 57
rect 1664 53 1670 54
rect 1674 53 1682 57
rect 1664 51 1682 53
rect 1607 49 1617 50
rect 1102 47 1117 48
rect 1106 43 1117 47
rect 1102 42 1117 43
rect 1119 47 1139 48
rect 1119 43 1135 47
rect 1119 42 1139 43
rect 1146 47 1156 48
rect 1146 43 1148 47
rect 1152 43 1156 47
rect 1146 42 1156 43
rect 1158 47 1177 48
rect 1158 43 1165 47
rect 1169 43 1177 47
rect 1158 42 1177 43
rect 1179 47 1187 48
rect 1179 43 1182 47
rect 1186 43 1187 47
rect 1179 42 1187 43
rect 1200 47 1210 48
rect 1200 43 1202 47
rect 1206 43 1210 47
rect 1200 42 1210 43
rect 1212 47 1231 48
rect 1212 43 1219 47
rect 1223 43 1231 47
rect 1212 42 1231 43
rect 1233 47 1241 48
rect 1233 43 1236 47
rect 1240 43 1241 47
rect 1233 42 1241 43
rect 1256 47 1266 48
rect 1256 43 1258 47
rect 1262 43 1266 47
rect 1256 42 1266 43
rect 1268 47 1287 48
rect 1268 43 1275 47
rect 1279 43 1287 47
rect 1268 42 1287 43
rect 1289 47 1297 48
rect 1289 43 1292 47
rect 1296 43 1297 47
rect 1289 42 1297 43
rect 1310 47 1320 48
rect 1310 43 1312 47
rect 1316 43 1320 47
rect 1310 42 1320 43
rect 1322 47 1341 48
rect 1322 43 1329 47
rect 1333 43 1341 47
rect 1322 42 1341 43
rect 1343 47 1351 48
rect 1343 43 1346 47
rect 1350 43 1351 47
rect 1343 42 1351 43
rect 1664 47 1682 49
rect 1664 43 1677 47
rect 1681 43 1682 47
rect 1664 41 1682 43
rect 1664 37 1682 39
rect 1655 31 1682 37
rect 1655 27 1656 31
rect 1660 27 1663 31
rect 1667 27 1682 31
rect 1655 25 1682 27
rect 1655 21 1682 23
rect 1655 18 1677 21
rect 1676 17 1677 18
rect 1681 17 1682 21
rect 1676 16 1682 17
rect 1512 -9 1518 -8
rect 1512 -10 1513 -9
rect 1505 -13 1513 -10
rect 1517 -10 1518 -9
rect 1517 -13 1523 -10
rect 1505 -15 1523 -13
rect 1505 -22 1523 -17
rect 1505 -27 1523 -24
rect 1505 -31 1506 -27
rect 1510 -31 1526 -27
rect 1505 -33 1526 -31
rect 1514 -35 1526 -33
rect 1514 -39 1526 -37
rect 1514 -43 1515 -39
rect 1519 -42 1526 -39
rect 1519 -43 1520 -42
rect 1514 -44 1520 -43
rect 1608 -2 1614 -1
rect 1608 -6 1609 -2
rect 1613 -3 1614 -2
rect 1613 -6 1635 -3
rect 1608 -8 1635 -6
rect 1608 -12 1635 -10
rect 1608 -16 1623 -12
rect 1627 -16 1630 -12
rect 1634 -16 1635 -12
rect 1608 -22 1635 -16
rect 1661 -17 1667 -16
rect 1661 -18 1662 -17
rect 1655 -21 1662 -18
rect 1666 -18 1667 -17
rect 1666 -21 1682 -18
rect 1608 -24 1626 -22
rect 1655 -23 1682 -21
rect 1608 -28 1626 -26
rect 1655 -27 1682 -25
rect 1608 -32 1609 -28
rect 1613 -32 1626 -28
rect 1608 -34 1626 -32
rect 1655 -30 1670 -27
rect 1664 -31 1670 -30
rect 1674 -31 1682 -27
rect 1664 -33 1682 -31
rect 1608 -38 1626 -36
rect 1608 -42 1616 -38
rect 1620 -39 1626 -38
rect 1620 -42 1635 -39
rect 1664 -37 1682 -35
rect 1664 -41 1677 -37
rect 1681 -41 1682 -37
rect 1608 -44 1635 -42
rect 1664 -43 1682 -41
rect 1608 -48 1635 -46
rect 1664 -47 1682 -45
rect 1608 -51 1624 -48
rect 1623 -52 1624 -51
rect 1628 -51 1635 -48
rect 1628 -52 1629 -51
rect 1623 -53 1629 -52
rect 1655 -53 1682 -47
rect 1655 -57 1656 -53
rect 1660 -57 1663 -53
rect 1667 -57 1682 -53
rect 1655 -59 1682 -57
rect 1655 -63 1682 -61
rect 1655 -66 1677 -63
rect 1676 -67 1677 -66
rect 1681 -67 1682 -63
rect 1676 -68 1682 -67
rect 1770 -26 1776 -25
rect 1770 -27 1771 -26
rect 1764 -30 1771 -27
rect 1775 -30 1776 -26
rect 1764 -32 1776 -30
rect 1764 -36 1776 -34
rect 1764 -38 1785 -36
rect 1764 -42 1780 -38
rect 1784 -42 1785 -38
rect 1767 -45 1785 -42
rect 1767 -52 1785 -47
rect 1767 -56 1785 -54
rect 1767 -59 1773 -56
rect 1772 -60 1773 -59
rect 1777 -59 1785 -56
rect 1777 -60 1778 -59
rect 1772 -61 1778 -60
rect 1032 -78 1063 -77
rect 146 -103 152 -96
rect 125 -111 132 -103
rect 125 -115 126 -111
rect 130 -115 132 -111
rect 125 -116 132 -115
rect 134 -104 142 -103
rect 134 -108 136 -104
rect 140 -108 142 -104
rect 134 -111 142 -108
rect 134 -115 136 -111
rect 140 -115 142 -111
rect 134 -116 142 -115
rect 144 -109 152 -103
rect 144 -113 146 -109
rect 150 -113 152 -109
rect 144 -114 152 -113
rect 154 -97 161 -96
rect 154 -101 156 -97
rect 160 -101 161 -97
rect 154 -104 161 -101
rect 233 -103 239 -96
rect 154 -108 156 -104
rect 160 -108 161 -104
rect 154 -109 161 -108
rect 154 -114 159 -109
rect 212 -111 219 -103
rect 144 -116 150 -114
rect 212 -115 213 -111
rect 217 -115 219 -111
rect 212 -116 219 -115
rect 221 -104 229 -103
rect 221 -108 223 -104
rect 227 -108 229 -104
rect 221 -111 229 -108
rect 221 -115 223 -111
rect 227 -115 229 -111
rect 221 -116 229 -115
rect 231 -109 239 -103
rect 231 -113 233 -109
rect 237 -113 239 -109
rect 231 -114 239 -113
rect 241 -97 248 -96
rect 241 -101 243 -97
rect 247 -101 248 -97
rect 241 -104 248 -101
rect 545 -95 552 -94
rect 326 -103 332 -96
rect 241 -108 243 -104
rect 247 -108 248 -104
rect 241 -109 248 -108
rect 241 -114 246 -109
rect 305 -111 312 -103
rect 231 -116 237 -114
rect 305 -115 306 -111
rect 310 -115 312 -111
rect 305 -116 312 -115
rect 314 -104 322 -103
rect 314 -108 316 -104
rect 320 -108 322 -104
rect 314 -111 322 -108
rect 314 -115 316 -111
rect 320 -115 322 -111
rect 314 -116 322 -115
rect 324 -109 332 -103
rect 324 -113 326 -109
rect 330 -113 332 -109
rect 324 -114 332 -113
rect 334 -97 341 -96
rect 334 -101 336 -97
rect 340 -101 341 -97
rect 334 -104 341 -101
rect 334 -108 336 -104
rect 340 -108 341 -104
rect 545 -99 546 -95
rect 550 -99 552 -95
rect 545 -102 552 -99
rect 545 -106 546 -102
rect 550 -106 552 -102
rect 545 -107 552 -106
rect 334 -109 341 -108
rect 334 -114 339 -109
rect 547 -112 552 -107
rect 554 -101 560 -94
rect 638 -95 645 -94
rect 638 -99 639 -95
rect 643 -99 645 -95
rect 554 -107 562 -101
rect 554 -111 556 -107
rect 560 -111 562 -107
rect 554 -112 562 -111
rect 324 -116 330 -114
rect 556 -114 562 -112
rect 564 -102 572 -101
rect 564 -106 566 -102
rect 570 -106 572 -102
rect 564 -109 572 -106
rect 564 -113 566 -109
rect 570 -113 572 -109
rect 564 -114 572 -113
rect 574 -109 581 -101
rect 638 -102 645 -99
rect 638 -106 639 -102
rect 643 -106 645 -102
rect 638 -107 645 -106
rect 574 -113 576 -109
rect 580 -113 581 -109
rect 640 -112 645 -107
rect 647 -101 653 -94
rect 725 -95 732 -94
rect 725 -99 726 -95
rect 730 -99 732 -95
rect 647 -107 655 -101
rect 647 -111 649 -107
rect 653 -111 655 -107
rect 647 -112 655 -111
rect 574 -114 581 -113
rect 649 -114 655 -112
rect 657 -102 665 -101
rect 657 -106 659 -102
rect 663 -106 665 -102
rect 657 -109 665 -106
rect 657 -113 659 -109
rect 663 -113 665 -109
rect 657 -114 665 -113
rect 667 -109 674 -101
rect 725 -102 732 -99
rect 725 -106 726 -102
rect 730 -106 732 -102
rect 725 -107 732 -106
rect 667 -113 669 -109
rect 673 -113 674 -109
rect 727 -112 732 -107
rect 734 -101 740 -94
rect 1032 -82 1037 -78
rect 1041 -82 1063 -78
rect 1032 -83 1063 -82
rect 1065 -82 1081 -77
rect 1087 -82 1100 -77
rect 1065 -83 1100 -82
rect 1120 -78 1135 -77
rect 1124 -82 1135 -78
rect 1120 -83 1135 -82
rect 1137 -78 1157 -77
rect 1137 -82 1153 -78
rect 1137 -83 1157 -82
rect 1164 -78 1174 -77
rect 1164 -82 1166 -78
rect 1170 -82 1174 -78
rect 1164 -83 1174 -82
rect 1176 -78 1195 -77
rect 1176 -82 1183 -78
rect 1187 -82 1195 -78
rect 1176 -83 1195 -82
rect 1197 -78 1205 -77
rect 1197 -82 1200 -78
rect 1204 -82 1205 -78
rect 1197 -83 1205 -82
rect 1218 -78 1228 -77
rect 1218 -82 1220 -78
rect 1224 -82 1228 -78
rect 1218 -83 1228 -82
rect 1230 -78 1249 -77
rect 1230 -82 1237 -78
rect 1241 -82 1249 -78
rect 1230 -83 1249 -82
rect 1251 -78 1259 -77
rect 1251 -82 1254 -78
rect 1258 -82 1259 -78
rect 1251 -83 1259 -82
rect 1274 -78 1284 -77
rect 1274 -82 1276 -78
rect 1280 -82 1284 -78
rect 1274 -83 1284 -82
rect 1286 -78 1305 -77
rect 1286 -82 1293 -78
rect 1297 -82 1305 -78
rect 1286 -83 1305 -82
rect 1307 -78 1315 -77
rect 1307 -82 1310 -78
rect 1314 -82 1315 -78
rect 1307 -83 1315 -82
rect 1328 -78 1338 -77
rect 1328 -82 1330 -78
rect 1334 -82 1338 -78
rect 1328 -83 1338 -82
rect 1340 -78 1359 -77
rect 1340 -82 1347 -78
rect 1351 -82 1359 -78
rect 1340 -83 1359 -82
rect 1361 -78 1369 -77
rect 1361 -82 1364 -78
rect 1368 -82 1369 -78
rect 1361 -83 1369 -82
rect 734 -107 742 -101
rect 734 -111 736 -107
rect 740 -111 742 -107
rect 734 -112 742 -111
rect 667 -114 674 -113
rect 736 -114 742 -112
rect 744 -102 752 -101
rect 744 -106 746 -102
rect 750 -106 752 -102
rect 744 -109 752 -106
rect 744 -113 746 -109
rect 750 -113 752 -109
rect 744 -114 752 -113
rect 754 -109 761 -101
rect 754 -113 756 -109
rect 760 -113 761 -109
rect 754 -114 761 -113
rect 1608 -86 1614 -85
rect 1608 -90 1609 -86
rect 1613 -87 1614 -86
rect 1613 -90 1635 -87
rect 1608 -92 1635 -90
rect 1608 -96 1635 -94
rect 1608 -100 1623 -96
rect 1627 -100 1630 -96
rect 1634 -100 1635 -96
rect 1608 -106 1635 -100
rect 1608 -108 1626 -106
rect 1608 -112 1626 -110
rect 1608 -116 1609 -112
rect 1613 -116 1626 -112
rect 1608 -118 1626 -116
rect 1673 -119 1683 -118
rect 1608 -122 1626 -120
rect 1608 -126 1616 -122
rect 1620 -123 1626 -122
rect 1620 -126 1635 -123
rect 1608 -128 1635 -126
rect 49 -164 54 -158
rect 47 -165 54 -164
rect 47 -169 48 -165
rect 52 -169 54 -165
rect 47 -170 54 -169
rect 56 -160 62 -158
rect 56 -165 64 -160
rect 56 -169 58 -165
rect 62 -169 64 -165
rect 56 -170 64 -169
rect 66 -165 74 -160
rect 66 -169 68 -165
rect 72 -169 74 -165
rect 66 -170 74 -169
rect 76 -161 83 -160
rect 76 -165 78 -161
rect 82 -165 83 -161
rect 135 -163 140 -142
rect 76 -170 83 -165
rect 133 -164 140 -163
rect 133 -168 134 -164
rect 138 -168 140 -164
rect 133 -169 140 -168
rect 142 -143 154 -142
rect 142 -147 144 -143
rect 148 -147 154 -143
rect 142 -150 154 -147
rect 142 -154 144 -150
rect 148 -151 154 -150
rect 171 -151 176 -142
rect 148 -154 156 -151
rect 142 -169 156 -154
rect 158 -164 166 -151
rect 158 -168 160 -164
rect 164 -168 166 -164
rect 158 -169 166 -168
rect 168 -157 176 -151
rect 168 -161 170 -157
rect 174 -161 176 -157
rect 168 -169 176 -161
rect 178 -148 183 -142
rect 178 -149 185 -148
rect 178 -153 180 -149
rect 184 -153 185 -149
rect 178 -154 185 -153
rect 178 -169 183 -154
rect 219 -163 224 -142
rect 217 -164 224 -163
rect 217 -168 218 -164
rect 222 -168 224 -164
rect 217 -169 224 -168
rect 226 -143 238 -142
rect 226 -147 228 -143
rect 232 -147 238 -143
rect 226 -150 238 -147
rect 226 -154 228 -150
rect 232 -151 238 -150
rect 255 -151 260 -142
rect 232 -154 240 -151
rect 226 -169 240 -154
rect 242 -164 250 -151
rect 242 -168 244 -164
rect 248 -168 250 -164
rect 242 -169 250 -168
rect 252 -157 260 -151
rect 252 -161 254 -157
rect 258 -161 260 -157
rect 252 -169 260 -161
rect 262 -148 267 -142
rect 262 -149 269 -148
rect 262 -153 264 -149
rect 268 -153 269 -149
rect 262 -154 269 -153
rect 262 -169 267 -154
rect 281 -164 286 -158
rect 279 -165 286 -164
rect 279 -169 280 -165
rect 284 -169 286 -165
rect 279 -170 286 -169
rect 288 -160 294 -158
rect 288 -165 296 -160
rect 288 -169 290 -165
rect 294 -169 296 -165
rect 288 -170 296 -169
rect 298 -165 306 -160
rect 298 -169 300 -165
rect 304 -169 306 -165
rect 298 -170 306 -169
rect 308 -161 315 -160
rect 308 -165 310 -161
rect 314 -165 315 -161
rect 378 -162 383 -156
rect 308 -170 315 -165
rect 376 -163 383 -162
rect 376 -167 377 -163
rect 381 -167 383 -163
rect 376 -168 383 -167
rect 385 -158 391 -156
rect 385 -163 393 -158
rect 385 -167 387 -163
rect 391 -167 393 -163
rect 385 -168 393 -167
rect 395 -163 403 -158
rect 395 -167 397 -163
rect 401 -167 403 -163
rect 395 -168 403 -167
rect 405 -159 412 -158
rect 405 -163 407 -159
rect 411 -163 412 -159
rect 464 -161 469 -140
rect 405 -168 412 -163
rect 462 -162 469 -161
rect 462 -166 463 -162
rect 467 -166 469 -162
rect 462 -167 469 -166
rect 471 -141 483 -140
rect 471 -145 473 -141
rect 477 -145 483 -141
rect 471 -148 483 -145
rect 471 -152 473 -148
rect 477 -149 483 -148
rect 500 -149 505 -140
rect 477 -152 485 -149
rect 471 -167 485 -152
rect 487 -162 495 -149
rect 487 -166 489 -162
rect 493 -166 495 -162
rect 487 -167 495 -166
rect 497 -155 505 -149
rect 497 -159 499 -155
rect 503 -159 505 -155
rect 497 -167 505 -159
rect 507 -146 512 -140
rect 507 -147 514 -146
rect 507 -151 509 -147
rect 513 -151 514 -147
rect 507 -152 514 -151
rect 507 -167 512 -152
rect 548 -161 553 -140
rect 546 -162 553 -161
rect 546 -166 547 -162
rect 551 -166 553 -162
rect 546 -167 553 -166
rect 555 -141 567 -140
rect 555 -145 557 -141
rect 561 -145 567 -141
rect 555 -148 567 -145
rect 555 -152 557 -148
rect 561 -149 567 -148
rect 584 -149 589 -140
rect 561 -152 569 -149
rect 555 -167 569 -152
rect 571 -162 579 -149
rect 571 -166 573 -162
rect 577 -166 579 -162
rect 571 -167 579 -166
rect 581 -155 589 -149
rect 581 -159 583 -155
rect 587 -159 589 -155
rect 581 -167 589 -159
rect 591 -146 596 -140
rect 591 -147 598 -146
rect 591 -151 593 -147
rect 597 -151 598 -147
rect 591 -152 598 -151
rect 591 -167 596 -152
rect 610 -162 615 -156
rect 608 -163 615 -162
rect 608 -167 609 -163
rect 613 -167 615 -163
rect 608 -168 615 -167
rect 617 -158 623 -156
rect 617 -163 625 -158
rect 617 -167 619 -163
rect 623 -167 625 -163
rect 617 -168 625 -167
rect 627 -163 635 -158
rect 627 -167 629 -163
rect 633 -167 635 -163
rect 627 -168 635 -167
rect 637 -159 644 -158
rect 705 -159 710 -153
rect 637 -163 639 -159
rect 643 -163 644 -159
rect 637 -168 644 -163
rect 703 -160 710 -159
rect 703 -164 704 -160
rect 708 -164 710 -160
rect 703 -165 710 -164
rect 712 -155 718 -153
rect 712 -160 720 -155
rect 712 -164 714 -160
rect 718 -164 720 -160
rect 712 -165 720 -164
rect 722 -160 730 -155
rect 722 -164 724 -160
rect 728 -164 730 -160
rect 722 -165 730 -164
rect 732 -156 739 -155
rect 732 -160 734 -156
rect 738 -160 739 -156
rect 791 -158 796 -137
rect 732 -165 739 -160
rect 789 -159 796 -158
rect 789 -163 790 -159
rect 794 -163 796 -159
rect 789 -164 796 -163
rect 798 -138 810 -137
rect 798 -142 800 -138
rect 804 -142 810 -138
rect 798 -145 810 -142
rect 798 -149 800 -145
rect 804 -146 810 -145
rect 827 -146 832 -137
rect 804 -149 812 -146
rect 798 -164 812 -149
rect 814 -159 822 -146
rect 814 -163 816 -159
rect 820 -163 822 -159
rect 814 -164 822 -163
rect 824 -152 832 -146
rect 824 -156 826 -152
rect 830 -156 832 -152
rect 824 -164 832 -156
rect 834 -143 839 -137
rect 834 -144 841 -143
rect 834 -148 836 -144
rect 840 -148 841 -144
rect 834 -149 841 -148
rect 834 -164 839 -149
rect 875 -158 880 -137
rect 873 -159 880 -158
rect 873 -163 874 -159
rect 878 -163 880 -159
rect 873 -164 880 -163
rect 882 -138 894 -137
rect 882 -142 884 -138
rect 888 -142 894 -138
rect 882 -145 894 -142
rect 882 -149 884 -145
rect 888 -146 894 -145
rect 911 -146 916 -137
rect 888 -149 896 -146
rect 882 -164 896 -149
rect 898 -159 906 -146
rect 898 -163 900 -159
rect 904 -163 906 -159
rect 898 -164 906 -163
rect 908 -152 916 -146
rect 908 -156 910 -152
rect 914 -156 916 -152
rect 908 -164 916 -156
rect 918 -143 923 -137
rect 1608 -132 1635 -130
rect 1608 -135 1624 -132
rect 1623 -136 1624 -135
rect 1628 -135 1635 -132
rect 1673 -123 1674 -119
rect 1678 -123 1683 -119
rect 1673 -125 1683 -123
rect 1673 -129 1683 -127
rect 1628 -136 1629 -135
rect 1623 -137 1629 -136
rect 1673 -133 1678 -129
rect 1682 -133 1683 -129
rect 1673 -135 1683 -133
rect 918 -144 925 -143
rect 918 -148 920 -144
rect 924 -148 925 -144
rect 918 -149 925 -148
rect 918 -164 923 -149
rect 937 -159 942 -153
rect 935 -160 942 -159
rect 935 -164 936 -160
rect 940 -164 942 -160
rect 935 -165 942 -164
rect 944 -155 950 -153
rect 944 -160 952 -155
rect 944 -164 946 -160
rect 950 -164 952 -160
rect 944 -165 952 -164
rect 954 -160 962 -155
rect 954 -164 956 -160
rect 960 -164 962 -160
rect 954 -165 962 -164
rect 964 -156 971 -155
rect 964 -160 966 -156
rect 970 -160 971 -156
rect 1607 -148 1613 -147
rect 1673 -139 1683 -137
rect 1671 -143 1678 -139
rect 1682 -143 1683 -139
rect 1671 -145 1683 -143
rect 1607 -152 1608 -148
rect 1612 -149 1613 -148
rect 1612 -152 1619 -149
rect 1607 -154 1619 -152
rect 1671 -149 1683 -147
rect 1671 -152 1678 -149
rect 1677 -153 1678 -152
rect 1682 -153 1683 -149
rect 964 -165 971 -160
rect 1607 -158 1619 -156
rect 1607 -162 1608 -158
rect 1612 -162 1619 -158
rect 1607 -164 1617 -162
rect 1677 -154 1683 -153
rect 1607 -168 1617 -166
rect 1607 -172 1608 -168
rect 1612 -172 1617 -168
rect 1607 -174 1617 -172
rect 1124 -177 1139 -176
rect 1128 -181 1139 -177
rect 1124 -182 1139 -181
rect 1141 -177 1161 -176
rect 1141 -181 1157 -177
rect 1141 -182 1161 -181
rect 1168 -177 1178 -176
rect 1168 -181 1170 -177
rect 1174 -181 1178 -177
rect 1168 -182 1178 -181
rect 1180 -177 1199 -176
rect 1180 -181 1187 -177
rect 1191 -181 1199 -177
rect 1180 -182 1199 -181
rect 1201 -177 1209 -176
rect 1201 -181 1204 -177
rect 1208 -181 1209 -177
rect 1201 -182 1209 -181
rect 1222 -177 1232 -176
rect 1222 -181 1224 -177
rect 1228 -181 1232 -177
rect 1222 -182 1232 -181
rect 1234 -177 1253 -176
rect 1234 -181 1241 -177
rect 1245 -181 1253 -177
rect 1234 -182 1253 -181
rect 1255 -177 1263 -176
rect 1255 -181 1258 -177
rect 1262 -181 1263 -177
rect 1255 -182 1263 -181
rect 1278 -177 1288 -176
rect 1278 -181 1280 -177
rect 1284 -181 1288 -177
rect 1278 -182 1288 -181
rect 1290 -177 1309 -176
rect 1290 -181 1297 -177
rect 1301 -181 1309 -177
rect 1290 -182 1309 -181
rect 1311 -177 1319 -176
rect 1311 -181 1314 -177
rect 1318 -181 1319 -177
rect 1311 -182 1319 -181
rect 1332 -177 1342 -176
rect 1332 -181 1334 -177
rect 1338 -181 1342 -177
rect 1332 -182 1342 -181
rect 1344 -177 1363 -176
rect 1344 -181 1351 -177
rect 1355 -181 1363 -177
rect 1344 -182 1363 -181
rect 1365 -177 1373 -176
rect 1365 -181 1368 -177
rect 1372 -181 1373 -177
rect 1365 -182 1373 -181
rect 1607 -178 1617 -176
rect 1607 -182 1612 -178
rect 1616 -182 1617 -178
rect 1607 -183 1617 -182
rect 159 -254 167 -251
rect 142 -259 147 -254
rect 140 -260 147 -259
rect 140 -264 141 -260
rect 145 -264 147 -260
rect 140 -265 147 -264
rect 142 -272 147 -265
rect 149 -272 154 -254
rect 156 -263 167 -254
rect 169 -257 174 -251
rect 1030 -223 1061 -222
rect 1030 -227 1035 -223
rect 1039 -227 1061 -223
rect 1030 -228 1061 -227
rect 1063 -227 1079 -222
rect 1085 -227 1098 -222
rect 1063 -228 1098 -227
rect 1118 -223 1133 -222
rect 1122 -227 1133 -223
rect 1118 -228 1133 -227
rect 1135 -223 1155 -222
rect 1135 -227 1151 -223
rect 1135 -228 1155 -227
rect 1162 -223 1172 -222
rect 1162 -227 1164 -223
rect 1168 -227 1172 -223
rect 1162 -228 1172 -227
rect 1174 -223 1193 -222
rect 1174 -227 1181 -223
rect 1185 -227 1193 -223
rect 1174 -228 1193 -227
rect 1195 -223 1203 -222
rect 1195 -227 1198 -223
rect 1202 -227 1203 -223
rect 1195 -228 1203 -227
rect 1216 -223 1226 -222
rect 1216 -227 1218 -223
rect 1222 -227 1226 -223
rect 1216 -228 1226 -227
rect 1228 -223 1247 -222
rect 1228 -227 1235 -223
rect 1239 -227 1247 -223
rect 1228 -228 1247 -227
rect 1249 -223 1257 -222
rect 1249 -227 1252 -223
rect 1256 -227 1257 -223
rect 1249 -228 1257 -227
rect 1272 -223 1282 -222
rect 1272 -227 1274 -223
rect 1278 -227 1282 -223
rect 1272 -228 1282 -227
rect 1284 -223 1303 -222
rect 1284 -227 1291 -223
rect 1295 -227 1303 -223
rect 1284 -228 1303 -227
rect 1305 -223 1313 -222
rect 1305 -227 1308 -223
rect 1312 -227 1313 -223
rect 1305 -228 1313 -227
rect 1326 -223 1336 -222
rect 1326 -227 1328 -223
rect 1332 -227 1336 -223
rect 1326 -228 1336 -227
rect 1338 -223 1357 -222
rect 1338 -227 1345 -223
rect 1349 -227 1357 -223
rect 1338 -228 1357 -227
rect 1359 -223 1367 -222
rect 1359 -227 1362 -223
rect 1366 -227 1367 -223
rect 1359 -228 1367 -227
rect 815 -249 823 -246
rect 488 -252 496 -249
rect 471 -257 476 -252
rect 169 -258 176 -257
rect 169 -262 171 -258
rect 175 -262 176 -258
rect 169 -263 176 -262
rect 469 -258 476 -257
rect 469 -262 470 -258
rect 474 -262 476 -258
rect 469 -263 476 -262
rect 156 -267 165 -263
rect 156 -271 159 -267
rect 163 -271 165 -267
rect 156 -272 165 -271
rect 471 -270 476 -263
rect 478 -270 483 -252
rect 485 -261 496 -252
rect 498 -255 503 -249
rect 798 -254 803 -249
rect 796 -255 803 -254
rect 498 -256 505 -255
rect 498 -260 500 -256
rect 504 -260 505 -256
rect 796 -259 797 -255
rect 801 -259 803 -255
rect 796 -260 803 -259
rect 498 -261 505 -260
rect 485 -265 494 -261
rect 485 -269 488 -265
rect 492 -269 494 -265
rect 798 -267 803 -260
rect 805 -267 810 -249
rect 812 -258 823 -249
rect 825 -252 830 -246
rect 825 -253 832 -252
rect 825 -257 827 -253
rect 831 -257 832 -253
rect 825 -258 832 -257
rect 812 -262 821 -258
rect 812 -266 815 -262
rect 819 -266 821 -262
rect 812 -267 821 -266
rect 485 -270 494 -269
rect 1665 -243 1675 -242
rect 1665 -247 1666 -243
rect 1670 -247 1675 -243
rect 1665 -249 1675 -247
rect 1665 -253 1675 -251
rect 1665 -257 1670 -253
rect 1674 -257 1675 -253
rect 1665 -259 1675 -257
rect 1410 -277 1415 -270
rect 1408 -278 1415 -277
rect 48 -310 53 -304
rect 46 -311 53 -310
rect 46 -315 47 -311
rect 51 -315 53 -311
rect 46 -316 53 -315
rect 55 -306 61 -304
rect 55 -311 63 -306
rect 55 -315 57 -311
rect 61 -315 63 -311
rect 55 -316 63 -315
rect 65 -311 73 -306
rect 65 -315 67 -311
rect 71 -315 73 -311
rect 65 -316 73 -315
rect 75 -307 82 -306
rect 75 -311 77 -307
rect 81 -311 82 -307
rect 134 -309 139 -288
rect 75 -316 82 -311
rect 132 -310 139 -309
rect 132 -314 133 -310
rect 137 -314 139 -310
rect 132 -315 139 -314
rect 141 -289 153 -288
rect 141 -293 143 -289
rect 147 -293 153 -289
rect 141 -296 153 -293
rect 141 -300 143 -296
rect 147 -297 153 -296
rect 170 -297 175 -288
rect 147 -300 155 -297
rect 141 -315 155 -300
rect 157 -310 165 -297
rect 157 -314 159 -310
rect 163 -314 165 -310
rect 157 -315 165 -314
rect 167 -303 175 -297
rect 167 -307 169 -303
rect 173 -307 175 -303
rect 167 -315 175 -307
rect 177 -294 182 -288
rect 177 -295 184 -294
rect 177 -299 179 -295
rect 183 -299 184 -295
rect 177 -300 184 -299
rect 177 -315 182 -300
rect 218 -309 223 -288
rect 216 -310 223 -309
rect 216 -314 217 -310
rect 221 -314 223 -310
rect 216 -315 223 -314
rect 225 -289 237 -288
rect 225 -293 227 -289
rect 231 -293 237 -289
rect 225 -296 237 -293
rect 225 -300 227 -296
rect 231 -297 237 -296
rect 254 -297 259 -288
rect 231 -300 239 -297
rect 225 -315 239 -300
rect 241 -310 249 -297
rect 241 -314 243 -310
rect 247 -314 249 -310
rect 241 -315 249 -314
rect 251 -303 259 -297
rect 251 -307 253 -303
rect 257 -307 259 -303
rect 251 -315 259 -307
rect 261 -294 266 -288
rect 261 -295 268 -294
rect 261 -299 263 -295
rect 267 -299 268 -295
rect 261 -300 268 -299
rect 261 -315 266 -300
rect 280 -310 285 -304
rect 278 -311 285 -310
rect 278 -315 279 -311
rect 283 -315 285 -311
rect 278 -316 285 -315
rect 287 -306 293 -304
rect 287 -311 295 -306
rect 287 -315 289 -311
rect 293 -315 295 -311
rect 287 -316 295 -315
rect 297 -311 305 -306
rect 297 -315 299 -311
rect 303 -315 305 -311
rect 297 -316 305 -315
rect 307 -307 314 -306
rect 307 -311 309 -307
rect 313 -311 314 -307
rect 377 -308 382 -302
rect 307 -316 314 -311
rect 375 -309 382 -308
rect 375 -313 376 -309
rect 380 -313 382 -309
rect 375 -314 382 -313
rect 384 -304 390 -302
rect 384 -309 392 -304
rect 384 -313 386 -309
rect 390 -313 392 -309
rect 384 -314 392 -313
rect 394 -309 402 -304
rect 394 -313 396 -309
rect 400 -313 402 -309
rect 394 -314 402 -313
rect 404 -305 411 -304
rect 404 -309 406 -305
rect 410 -309 411 -305
rect 463 -307 468 -286
rect 404 -314 411 -309
rect 461 -308 468 -307
rect 461 -312 462 -308
rect 466 -312 468 -308
rect 461 -313 468 -312
rect 470 -287 482 -286
rect 470 -291 472 -287
rect 476 -291 482 -287
rect 470 -294 482 -291
rect 470 -298 472 -294
rect 476 -295 482 -294
rect 499 -295 504 -286
rect 476 -298 484 -295
rect 470 -313 484 -298
rect 486 -308 494 -295
rect 486 -312 488 -308
rect 492 -312 494 -308
rect 486 -313 494 -312
rect 496 -301 504 -295
rect 496 -305 498 -301
rect 502 -305 504 -301
rect 496 -313 504 -305
rect 506 -292 511 -286
rect 506 -293 513 -292
rect 506 -297 508 -293
rect 512 -297 513 -293
rect 506 -298 513 -297
rect 506 -313 511 -298
rect 547 -307 552 -286
rect 545 -308 552 -307
rect 545 -312 546 -308
rect 550 -312 552 -308
rect 545 -313 552 -312
rect 554 -287 566 -286
rect 554 -291 556 -287
rect 560 -291 566 -287
rect 554 -294 566 -291
rect 554 -298 556 -294
rect 560 -295 566 -294
rect 583 -295 588 -286
rect 560 -298 568 -295
rect 554 -313 568 -298
rect 570 -308 578 -295
rect 570 -312 572 -308
rect 576 -312 578 -308
rect 570 -313 578 -312
rect 580 -301 588 -295
rect 580 -305 582 -301
rect 586 -305 588 -301
rect 580 -313 588 -305
rect 590 -292 595 -286
rect 590 -293 597 -292
rect 590 -297 592 -293
rect 596 -297 597 -293
rect 590 -298 597 -297
rect 590 -313 595 -298
rect 609 -308 614 -302
rect 607 -309 614 -308
rect 607 -313 608 -309
rect 612 -313 614 -309
rect 607 -314 614 -313
rect 616 -304 622 -302
rect 616 -309 624 -304
rect 616 -313 618 -309
rect 622 -313 624 -309
rect 616 -314 624 -313
rect 626 -309 634 -304
rect 626 -313 628 -309
rect 632 -313 634 -309
rect 626 -314 634 -313
rect 636 -305 643 -304
rect 704 -305 709 -299
rect 636 -309 638 -305
rect 642 -309 643 -305
rect 636 -314 643 -309
rect 702 -306 709 -305
rect 702 -310 703 -306
rect 707 -310 709 -306
rect 702 -311 709 -310
rect 711 -301 717 -299
rect 711 -306 719 -301
rect 711 -310 713 -306
rect 717 -310 719 -306
rect 711 -311 719 -310
rect 721 -306 729 -301
rect 721 -310 723 -306
rect 727 -310 729 -306
rect 721 -311 729 -310
rect 731 -302 738 -301
rect 731 -306 733 -302
rect 737 -306 738 -302
rect 790 -304 795 -283
rect 731 -311 738 -306
rect 788 -305 795 -304
rect 788 -309 789 -305
rect 793 -309 795 -305
rect 788 -310 795 -309
rect 797 -284 809 -283
rect 797 -288 799 -284
rect 803 -288 809 -284
rect 797 -291 809 -288
rect 797 -295 799 -291
rect 803 -292 809 -291
rect 826 -292 831 -283
rect 803 -295 811 -292
rect 797 -310 811 -295
rect 813 -305 821 -292
rect 813 -309 815 -305
rect 819 -309 821 -305
rect 813 -310 821 -309
rect 823 -298 831 -292
rect 823 -302 825 -298
rect 829 -302 831 -298
rect 823 -310 831 -302
rect 833 -289 838 -283
rect 833 -290 840 -289
rect 833 -294 835 -290
rect 839 -294 840 -290
rect 833 -295 840 -294
rect 833 -310 838 -295
rect 874 -304 879 -283
rect 872 -305 879 -304
rect 872 -309 873 -305
rect 877 -309 879 -305
rect 872 -310 879 -309
rect 881 -284 893 -283
rect 881 -288 883 -284
rect 887 -288 893 -284
rect 881 -291 893 -288
rect 881 -295 883 -291
rect 887 -292 893 -291
rect 910 -292 915 -283
rect 887 -295 895 -292
rect 881 -310 895 -295
rect 897 -305 905 -292
rect 897 -309 899 -305
rect 903 -309 905 -305
rect 897 -310 905 -309
rect 907 -298 915 -292
rect 907 -302 909 -298
rect 913 -302 915 -298
rect 907 -310 915 -302
rect 917 -289 922 -283
rect 1408 -282 1409 -278
rect 1413 -282 1415 -278
rect 1408 -283 1415 -282
rect 917 -290 924 -289
rect 917 -294 919 -290
rect 923 -294 924 -290
rect 917 -295 924 -294
rect 917 -310 922 -295
rect 936 -305 941 -299
rect 934 -306 941 -305
rect 934 -310 935 -306
rect 939 -310 941 -306
rect 934 -311 941 -310
rect 943 -301 949 -299
rect 943 -306 951 -301
rect 943 -310 945 -306
rect 949 -310 951 -306
rect 943 -311 951 -310
rect 953 -306 961 -301
rect 953 -310 955 -306
rect 959 -310 961 -306
rect 953 -311 961 -310
rect 963 -302 970 -301
rect 963 -306 965 -302
rect 969 -306 970 -302
rect 1410 -287 1415 -283
rect 1417 -287 1427 -270
rect 1419 -296 1427 -287
rect 1419 -300 1420 -296
rect 1424 -298 1427 -296
rect 1429 -278 1434 -270
rect 1665 -263 1675 -261
rect 1663 -267 1670 -263
rect 1674 -267 1675 -263
rect 1663 -269 1675 -267
rect 1663 -273 1675 -271
rect 1663 -276 1670 -273
rect 1669 -277 1670 -276
rect 1674 -277 1675 -273
rect 1669 -278 1675 -277
rect 1429 -279 1436 -278
rect 1429 -283 1431 -279
rect 1435 -283 1436 -279
rect 1429 -286 1436 -283
rect 1429 -290 1431 -286
rect 1435 -290 1436 -286
rect 1653 -289 1659 -288
rect 1653 -290 1654 -289
rect 1429 -291 1436 -290
rect 1429 -298 1434 -291
rect 1647 -293 1654 -290
rect 1658 -290 1659 -289
rect 1658 -293 1674 -290
rect 1647 -295 1674 -293
rect 1424 -300 1425 -298
rect 1419 -301 1425 -300
rect 1647 -299 1674 -297
rect 1647 -302 1662 -299
rect 1656 -303 1662 -302
rect 1666 -303 1674 -299
rect 1656 -305 1674 -303
rect 963 -311 970 -306
rect 1656 -309 1674 -307
rect 1656 -313 1669 -309
rect 1673 -313 1674 -309
rect 1656 -315 1674 -313
rect 1656 -319 1674 -317
rect 1122 -322 1137 -321
rect 1126 -326 1137 -322
rect 1122 -327 1137 -326
rect 1139 -322 1159 -321
rect 1139 -326 1155 -322
rect 1139 -327 1159 -326
rect 1166 -322 1176 -321
rect 1166 -326 1168 -322
rect 1172 -326 1176 -322
rect 1166 -327 1176 -326
rect 1178 -322 1197 -321
rect 1178 -326 1185 -322
rect 1189 -326 1197 -322
rect 1178 -327 1197 -326
rect 1199 -322 1207 -321
rect 1199 -326 1202 -322
rect 1206 -326 1207 -322
rect 1199 -327 1207 -326
rect 1220 -322 1230 -321
rect 1220 -326 1222 -322
rect 1226 -326 1230 -322
rect 1220 -327 1230 -326
rect 1232 -322 1251 -321
rect 1232 -326 1239 -322
rect 1243 -326 1251 -322
rect 1232 -327 1251 -326
rect 1253 -322 1261 -321
rect 1253 -326 1256 -322
rect 1260 -326 1261 -322
rect 1253 -327 1261 -326
rect 1276 -322 1286 -321
rect 1276 -326 1278 -322
rect 1282 -326 1286 -322
rect 1276 -327 1286 -326
rect 1288 -322 1307 -321
rect 1288 -326 1295 -322
rect 1299 -326 1307 -322
rect 1288 -327 1307 -326
rect 1309 -322 1317 -321
rect 1309 -326 1312 -322
rect 1316 -326 1317 -322
rect 1309 -327 1317 -326
rect 1330 -322 1340 -321
rect 1330 -326 1332 -322
rect 1336 -326 1340 -322
rect 1330 -327 1340 -326
rect 1342 -322 1361 -321
rect 1342 -326 1349 -322
rect 1353 -326 1361 -322
rect 1342 -327 1361 -326
rect 1363 -322 1371 -321
rect 1363 -326 1366 -322
rect 1370 -326 1371 -322
rect 1363 -327 1371 -326
rect 1647 -325 1674 -319
rect 1421 -329 1427 -328
rect 1421 -333 1422 -329
rect 1426 -331 1427 -329
rect 1647 -329 1648 -325
rect 1652 -329 1655 -325
rect 1659 -329 1674 -325
rect 1647 -331 1674 -329
rect 1426 -333 1429 -331
rect 1421 -342 1429 -333
rect 1412 -346 1417 -342
rect 1410 -347 1417 -346
rect 1410 -351 1411 -347
rect 1415 -351 1417 -347
rect 1410 -352 1417 -351
rect 1031 -365 1062 -364
rect 158 -400 166 -397
rect 141 -405 146 -400
rect 139 -406 146 -405
rect 139 -410 140 -406
rect 144 -410 146 -406
rect 139 -411 146 -410
rect 141 -418 146 -411
rect 148 -418 153 -400
rect 155 -409 166 -400
rect 168 -403 173 -397
rect 1031 -369 1036 -365
rect 1040 -369 1062 -365
rect 1031 -370 1062 -369
rect 1064 -369 1080 -364
rect 1412 -359 1417 -352
rect 1419 -359 1429 -342
rect 1431 -338 1436 -331
rect 1647 -335 1674 -333
rect 1647 -338 1669 -335
rect 1431 -339 1438 -338
rect 1431 -343 1433 -339
rect 1437 -343 1438 -339
rect 1668 -339 1669 -338
rect 1673 -339 1674 -335
rect 1668 -340 1674 -339
rect 1431 -346 1438 -343
rect 1431 -350 1433 -346
rect 1437 -350 1438 -346
rect 1431 -351 1438 -350
rect 1431 -359 1436 -351
rect 1086 -369 1099 -364
rect 1064 -370 1099 -369
rect 1119 -365 1134 -364
rect 1123 -369 1134 -365
rect 1119 -370 1134 -369
rect 1136 -365 1156 -364
rect 1136 -369 1152 -365
rect 1136 -370 1156 -369
rect 1163 -365 1173 -364
rect 1163 -369 1165 -365
rect 1169 -369 1173 -365
rect 1163 -370 1173 -369
rect 1175 -365 1194 -364
rect 1175 -369 1182 -365
rect 1186 -369 1194 -365
rect 1175 -370 1194 -369
rect 1196 -365 1204 -364
rect 1196 -369 1199 -365
rect 1203 -369 1204 -365
rect 1196 -370 1204 -369
rect 1217 -365 1227 -364
rect 1217 -369 1219 -365
rect 1223 -369 1227 -365
rect 1217 -370 1227 -369
rect 1229 -365 1248 -364
rect 1229 -369 1236 -365
rect 1240 -369 1248 -365
rect 1229 -370 1248 -369
rect 1250 -365 1258 -364
rect 1250 -369 1253 -365
rect 1257 -369 1258 -365
rect 1250 -370 1258 -369
rect 1273 -365 1283 -364
rect 1273 -369 1275 -365
rect 1279 -369 1283 -365
rect 1273 -370 1283 -369
rect 1285 -365 1304 -364
rect 1285 -369 1292 -365
rect 1296 -369 1304 -365
rect 1285 -370 1304 -369
rect 1306 -365 1314 -364
rect 1306 -369 1309 -365
rect 1313 -369 1314 -365
rect 1306 -370 1314 -369
rect 1327 -365 1337 -364
rect 1327 -369 1329 -365
rect 1333 -369 1337 -365
rect 1327 -370 1337 -369
rect 1339 -365 1358 -364
rect 1339 -369 1346 -365
rect 1350 -369 1358 -365
rect 1339 -370 1358 -369
rect 1360 -365 1368 -364
rect 1360 -369 1363 -365
rect 1367 -369 1368 -365
rect 1360 -370 1368 -369
rect 814 -395 822 -392
rect 487 -398 495 -395
rect 470 -403 475 -398
rect 168 -404 175 -403
rect 168 -408 170 -404
rect 174 -408 175 -404
rect 168 -409 175 -408
rect 468 -404 475 -403
rect 468 -408 469 -404
rect 473 -408 475 -404
rect 468 -409 475 -408
rect 155 -413 164 -409
rect 155 -417 158 -413
rect 162 -417 164 -413
rect 155 -418 164 -417
rect 470 -416 475 -409
rect 477 -416 482 -398
rect 484 -407 495 -398
rect 497 -401 502 -395
rect 797 -400 802 -395
rect 795 -401 802 -400
rect 497 -402 504 -401
rect 497 -406 499 -402
rect 503 -406 504 -402
rect 795 -405 796 -401
rect 800 -405 802 -401
rect 795 -406 802 -405
rect 497 -407 504 -406
rect 484 -411 493 -407
rect 484 -415 487 -411
rect 491 -415 493 -411
rect 797 -413 802 -406
rect 804 -413 809 -395
rect 811 -404 822 -395
rect 824 -398 829 -392
rect 824 -399 831 -398
rect 824 -403 826 -399
rect 830 -403 831 -399
rect 824 -404 831 -403
rect 811 -408 820 -404
rect 1653 -373 1659 -372
rect 1653 -374 1654 -373
rect 1647 -377 1654 -374
rect 1658 -374 1659 -373
rect 1658 -377 1674 -374
rect 1647 -379 1674 -377
rect 1647 -383 1674 -381
rect 811 -412 814 -408
rect 818 -412 820 -408
rect 1647 -386 1662 -383
rect 1656 -387 1662 -386
rect 1666 -387 1674 -383
rect 1656 -389 1674 -387
rect 1656 -393 1674 -391
rect 1656 -397 1669 -393
rect 1673 -397 1674 -393
rect 1656 -399 1674 -397
rect 1656 -403 1674 -401
rect 1647 -409 1674 -403
rect 811 -413 820 -412
rect 484 -416 493 -415
rect 1647 -413 1648 -409
rect 1652 -413 1655 -409
rect 1659 -413 1674 -409
rect 1647 -415 1674 -413
rect 351 -445 357 -443
rect 342 -450 347 -445
rect 340 -451 347 -450
rect 340 -455 341 -451
rect 345 -455 347 -451
rect 340 -458 347 -455
rect 340 -462 341 -458
rect 345 -462 347 -458
rect 340 -463 347 -462
rect 349 -446 357 -445
rect 349 -450 351 -446
rect 355 -450 357 -446
rect 349 -456 357 -450
rect 359 -444 367 -443
rect 359 -448 361 -444
rect 365 -448 367 -444
rect 359 -451 367 -448
rect 359 -455 361 -451
rect 365 -455 367 -451
rect 359 -456 367 -455
rect 369 -444 376 -443
rect 369 -448 371 -444
rect 375 -448 376 -444
rect 444 -445 450 -443
rect 369 -456 376 -448
rect 435 -450 440 -445
rect 433 -451 440 -450
rect 433 -455 434 -451
rect 438 -455 440 -451
rect 349 -463 355 -456
rect 433 -458 440 -455
rect 433 -462 434 -458
rect 438 -462 440 -458
rect 433 -463 440 -462
rect 442 -446 450 -445
rect 442 -450 444 -446
rect 448 -450 450 -446
rect 442 -456 450 -450
rect 452 -444 460 -443
rect 452 -448 454 -444
rect 458 -448 460 -444
rect 452 -451 460 -448
rect 452 -455 454 -451
rect 458 -455 460 -451
rect 452 -456 460 -455
rect 462 -444 469 -443
rect 462 -448 464 -444
rect 468 -448 469 -444
rect 531 -445 537 -443
rect 462 -456 469 -448
rect 522 -450 527 -445
rect 520 -451 527 -450
rect 520 -455 521 -451
rect 525 -455 527 -451
rect 442 -463 448 -456
rect 520 -458 527 -455
rect 520 -462 521 -458
rect 525 -462 527 -458
rect 520 -463 527 -462
rect 529 -446 537 -445
rect 529 -450 531 -446
rect 535 -450 537 -446
rect 529 -456 537 -450
rect 539 -444 547 -443
rect 539 -448 541 -444
rect 545 -448 547 -444
rect 539 -451 547 -448
rect 539 -455 541 -451
rect 545 -455 547 -451
rect 539 -456 547 -455
rect 549 -444 556 -443
rect 549 -448 551 -444
rect 555 -448 556 -444
rect 1647 -419 1674 -417
rect 1647 -422 1669 -419
rect 1668 -423 1669 -422
rect 1673 -423 1674 -419
rect 1668 -424 1674 -423
rect 1762 -382 1768 -381
rect 1762 -383 1763 -382
rect 1756 -386 1763 -383
rect 1767 -386 1768 -382
rect 1756 -388 1768 -386
rect 1756 -392 1768 -390
rect 1756 -394 1777 -392
rect 1756 -398 1772 -394
rect 1776 -398 1777 -394
rect 1759 -401 1777 -398
rect 1759 -408 1777 -403
rect 1759 -412 1777 -410
rect 1759 -415 1765 -412
rect 1764 -416 1765 -415
rect 1769 -415 1777 -412
rect 1769 -416 1770 -415
rect 1764 -417 1770 -416
rect 1751 -430 1768 -429
rect 1751 -434 1752 -430
rect 1756 -434 1759 -430
rect 1763 -431 1768 -430
rect 1763 -434 1776 -431
rect 1751 -436 1776 -434
rect 1751 -441 1776 -438
rect 549 -456 556 -448
rect 529 -463 535 -456
rect 1414 -456 1419 -449
rect 1412 -457 1419 -456
rect 1412 -461 1413 -457
rect 1417 -461 1419 -457
rect 1412 -462 1419 -461
rect 1123 -464 1138 -463
rect 1127 -468 1138 -464
rect 1123 -469 1138 -468
rect 1140 -464 1160 -463
rect 1140 -468 1156 -464
rect 1140 -469 1160 -468
rect 1167 -464 1177 -463
rect 1167 -468 1169 -464
rect 1173 -468 1177 -464
rect 1167 -469 1177 -468
rect 1179 -464 1198 -463
rect 1179 -468 1186 -464
rect 1190 -468 1198 -464
rect 1179 -469 1198 -468
rect 1200 -464 1208 -463
rect 1200 -468 1203 -464
rect 1207 -468 1208 -464
rect 1200 -469 1208 -468
rect 1221 -464 1231 -463
rect 1221 -468 1223 -464
rect 1227 -468 1231 -464
rect 1221 -469 1231 -468
rect 1233 -464 1252 -463
rect 1233 -468 1240 -464
rect 1244 -468 1252 -464
rect 1233 -469 1252 -468
rect 1254 -464 1262 -463
rect 1254 -468 1257 -464
rect 1261 -468 1262 -464
rect 1254 -469 1262 -468
rect 1277 -464 1287 -463
rect 1277 -468 1279 -464
rect 1283 -468 1287 -464
rect 1277 -469 1287 -468
rect 1289 -464 1308 -463
rect 1289 -468 1296 -464
rect 1300 -468 1308 -464
rect 1289 -469 1308 -468
rect 1310 -464 1318 -463
rect 1310 -468 1313 -464
rect 1317 -468 1318 -464
rect 1310 -469 1318 -468
rect 1331 -464 1341 -463
rect 1331 -468 1333 -464
rect 1337 -468 1341 -464
rect 1331 -469 1341 -468
rect 1343 -464 1362 -463
rect 1343 -468 1350 -464
rect 1354 -468 1362 -464
rect 1343 -469 1362 -468
rect 1364 -464 1372 -463
rect 1364 -468 1367 -464
rect 1371 -468 1372 -464
rect 1414 -466 1419 -462
rect 1421 -466 1431 -449
rect 1364 -469 1372 -468
rect 1423 -475 1431 -466
rect 1423 -479 1424 -475
rect 1428 -477 1431 -475
rect 1433 -457 1438 -449
rect 1751 -445 1772 -441
rect 1751 -447 1776 -445
rect 1751 -449 1764 -447
rect 1751 -453 1764 -451
rect 1751 -454 1752 -453
rect 1433 -458 1440 -457
rect 1433 -462 1435 -458
rect 1439 -462 1440 -458
rect 1433 -465 1440 -462
rect 1433 -469 1435 -465
rect 1439 -469 1440 -465
rect 1748 -457 1752 -454
rect 1756 -454 1764 -453
rect 1756 -457 1773 -454
rect 1748 -459 1773 -457
rect 1748 -466 1773 -461
rect 1433 -470 1440 -469
rect 1433 -477 1438 -470
rect 1665 -475 1675 -474
rect 1428 -479 1429 -477
rect 1423 -480 1429 -479
rect 1665 -479 1666 -475
rect 1670 -479 1675 -475
rect 1665 -481 1675 -479
rect 1665 -485 1675 -483
rect 1665 -489 1670 -485
rect 1674 -489 1675 -485
rect 1748 -470 1773 -468
rect 1748 -476 1776 -470
rect 1748 -480 1764 -476
rect 1768 -480 1771 -476
rect 1775 -480 1776 -476
rect 1748 -484 1776 -480
rect 1748 -488 1776 -486
rect 1665 -491 1675 -489
rect 1748 -492 1756 -488
rect 1760 -492 1763 -488
rect 1767 -492 1776 -488
rect 1665 -495 1675 -493
rect 1663 -499 1670 -495
rect 1674 -499 1675 -495
rect 1663 -501 1675 -499
rect 1748 -494 1776 -492
rect 1748 -498 1776 -496
rect 1748 -502 1764 -498
rect 1768 -502 1771 -498
rect 1775 -502 1776 -498
rect 1663 -505 1675 -503
rect 1663 -508 1670 -505
rect 1669 -509 1670 -508
rect 1674 -509 1675 -505
rect 1669 -510 1675 -509
rect 1748 -504 1776 -502
rect 1748 -508 1776 -506
rect 1748 -512 1749 -508
rect 1753 -512 1756 -508
rect 1760 -511 1776 -508
rect 1760 -512 1761 -511
rect 1748 -513 1761 -512
<< metal1 >>
rect 1496 479 1520 480
rect 1496 478 1649 479
rect 1496 475 1655 478
rect 33 458 474 462
rect 33 436 37 458
rect 516 456 778 460
rect 115 449 116 452
rect 516 454 520 456
rect 467 451 520 454
rect 331 449 457 450
rect 530 449 574 451
rect 115 448 457 449
rect 110 447 457 448
rect 524 448 574 449
rect 623 448 667 451
rect 710 450 754 451
rect 710 448 762 450
rect 524 447 762 448
rect 110 445 536 447
rect 110 441 134 445
rect 138 441 144 445
rect 148 441 221 445
rect 225 441 231 445
rect 235 441 314 445
rect 318 441 324 445
rect 328 444 536 445
rect 328 441 334 444
rect 530 443 536 444
rect 540 443 546 447
rect 550 444 629 447
rect 550 443 574 444
rect 623 443 629 444
rect 633 443 639 447
rect 643 444 716 447
rect 643 443 667 444
rect 710 443 716 444
rect 720 443 726 447
rect 730 444 762 447
rect 730 443 754 444
rect 774 441 778 456
rect 951 452 1366 455
rect 951 451 1002 452
rect 994 441 999 444
rect 467 436 498 440
rect 114 431 115 435
rect 119 431 134 435
rect 114 424 126 428
rect 121 419 126 424
rect 130 427 134 431
rect 138 433 150 436
rect 138 430 145 433
rect 149 429 150 433
rect 201 431 202 435
rect 206 431 221 435
rect 145 428 150 429
rect 130 423 142 427
rect 138 419 142 423
rect 121 415 128 419
rect 132 415 135 419
rect 114 402 118 411
rect 122 407 127 411
rect 138 404 142 415
rect 146 414 150 428
rect 202 424 213 428
rect 208 419 213 424
rect 217 427 221 431
rect 225 433 237 436
rect 225 430 232 433
rect 236 429 237 433
rect 294 431 295 435
rect 299 431 314 435
rect 232 428 237 429
rect 217 423 229 427
rect 225 419 229 423
rect 208 415 215 419
rect 219 415 222 419
rect 146 411 175 414
rect 146 410 150 411
rect 107 398 118 402
rect 125 402 142 404
rect 129 400 142 402
rect 145 409 150 410
rect 149 405 150 409
rect 145 402 150 405
rect 125 395 129 398
rect 149 398 150 402
rect 145 397 150 398
rect 114 391 115 395
rect 119 391 120 395
rect 114 385 120 391
rect 125 390 129 391
rect 134 393 135 397
rect 139 393 140 397
rect 134 385 140 393
rect 110 381 144 385
rect 148 381 154 385
rect 110 377 154 381
rect 111 370 115 377
rect 171 375 175 411
rect 201 401 205 411
rect 209 407 214 411
rect 225 404 229 415
rect 233 410 237 428
rect 295 424 306 428
rect 301 419 306 424
rect 310 427 314 431
rect 318 433 330 436
rect 534 435 546 438
rect 318 430 325 433
rect 329 429 330 433
rect 343 429 515 433
rect 520 429 521 433
rect 534 431 535 435
rect 539 432 546 435
rect 550 433 565 437
rect 569 433 570 437
rect 627 435 639 438
rect 534 430 539 431
rect 325 428 330 429
rect 310 423 322 427
rect 318 419 322 423
rect 301 415 308 419
rect 312 415 315 419
rect 198 398 205 401
rect 212 402 229 404
rect 216 400 229 402
rect 232 409 237 410
rect 236 405 237 409
rect 232 402 237 405
rect 212 395 216 398
rect 236 400 237 402
rect 236 398 243 400
rect 232 397 243 398
rect 294 401 298 411
rect 302 407 307 411
rect 318 404 322 415
rect 326 421 330 428
rect 534 423 538 430
rect 550 429 554 433
rect 627 431 628 435
rect 632 432 639 435
rect 643 433 658 437
rect 662 433 663 437
rect 714 435 726 438
rect 774 437 980 441
rect 627 430 632 431
rect 326 417 412 421
rect 478 419 538 423
rect 326 410 330 417
rect 534 412 538 419
rect 542 425 554 429
rect 558 427 569 430
rect 542 421 546 425
rect 558 421 563 427
rect 549 417 552 421
rect 556 417 563 421
rect 627 419 631 430
rect 643 429 647 433
rect 714 431 715 435
rect 719 432 726 435
rect 730 433 745 437
rect 749 433 750 437
rect 714 430 719 431
rect 534 411 539 412
rect 291 398 298 401
rect 305 402 322 404
rect 309 400 322 402
rect 325 409 330 410
rect 329 405 330 409
rect 343 407 516 410
rect 534 407 535 411
rect 325 402 330 405
rect 201 391 202 395
rect 206 391 207 395
rect 201 385 207 391
rect 212 390 216 391
rect 221 393 222 397
rect 226 393 227 397
rect 305 395 309 398
rect 329 398 330 402
rect 534 404 539 407
rect 534 400 535 404
rect 542 406 546 417
rect 604 416 631 419
rect 557 409 562 413
rect 542 404 559 406
rect 542 402 555 404
rect 534 399 539 400
rect 566 403 570 413
rect 604 404 608 416
rect 566 400 573 403
rect 325 397 330 398
rect 221 385 227 393
rect 294 391 295 395
rect 299 391 300 395
rect 294 385 300 391
rect 305 390 309 391
rect 314 393 315 397
rect 319 393 320 397
rect 544 395 545 399
rect 549 395 550 399
rect 314 385 320 393
rect 343 389 517 392
rect 544 387 550 395
rect 555 397 559 400
rect 627 412 631 416
rect 635 425 647 429
rect 651 429 665 430
rect 651 427 662 429
rect 635 421 639 425
rect 651 421 656 427
rect 642 417 645 421
rect 649 417 656 421
rect 627 411 632 412
rect 627 407 628 411
rect 627 404 632 407
rect 627 400 628 404
rect 635 406 639 417
rect 714 416 718 430
rect 730 429 734 433
rect 650 409 655 413
rect 635 404 652 406
rect 635 402 648 404
rect 627 399 632 400
rect 659 403 663 413
rect 692 412 718 416
rect 722 425 734 429
rect 738 429 752 430
rect 994 429 997 441
rect 1016 433 1019 452
rect 1029 441 1083 444
rect 1061 435 1065 437
rect 738 427 749 429
rect 722 421 726 425
rect 738 421 743 427
rect 753 425 998 429
rect 729 417 732 421
rect 736 417 743 421
rect 1061 418 1065 429
rect 1080 426 1083 441
rect 1099 433 1102 452
rect 1162 433 1165 452
rect 1172 447 1175 452
rect 1216 433 1219 452
rect 1226 447 1229 452
rect 1272 433 1275 452
rect 1282 447 1285 452
rect 1326 433 1329 452
rect 1336 447 1339 452
rect 1080 423 1130 426
rect 659 400 666 403
rect 678 402 679 406
rect 555 392 559 393
rect 564 393 565 397
rect 569 393 570 397
rect 564 387 570 393
rect 637 395 638 399
rect 642 395 643 399
rect 637 387 643 395
rect 648 397 652 400
rect 648 392 652 393
rect 657 393 658 397
rect 662 393 663 397
rect 657 387 663 393
rect 197 381 231 385
rect 235 381 241 385
rect 197 380 241 381
rect 290 381 324 385
rect 328 381 334 385
rect 197 377 224 380
rect 290 377 334 381
rect 530 383 536 387
rect 540 383 574 387
rect 623 383 629 387
rect 633 383 667 387
rect 530 379 574 383
rect 199 370 203 377
rect 236 373 269 376
rect 290 370 294 377
rect 566 375 570 379
rect 585 378 615 381
rect 623 379 667 383
rect 678 382 682 402
rect 524 374 628 375
rect 524 372 650 374
rect 659 372 663 379
rect 692 381 696 412
rect 714 411 719 412
rect 714 407 715 411
rect 702 382 706 402
rect 714 404 719 407
rect 714 400 715 404
rect 722 406 726 417
rect 737 409 742 413
rect 722 404 739 406
rect 722 402 735 404
rect 714 399 719 400
rect 746 404 750 413
rect 1044 414 1047 417
rect 1061 408 1064 418
rect 1116 413 1119 416
rect 746 400 754 404
rect 724 395 725 399
rect 729 395 730 399
rect 724 387 730 395
rect 735 397 739 400
rect 735 392 739 393
rect 744 393 745 397
rect 749 393 750 397
rect 744 387 750 393
rect 710 383 716 387
rect 720 383 754 387
rect 710 379 754 383
rect 748 372 752 379
rect 945 375 949 408
rect 1061 404 1062 408
rect 1061 396 1064 404
rect 1126 403 1130 423
rect 1133 407 1136 429
rect 1146 424 1149 429
rect 1179 424 1182 429
rect 1146 421 1182 424
rect 1148 413 1150 416
rect 1162 414 1166 416
rect 1170 414 1171 416
rect 1162 413 1171 414
rect 1133 403 1134 407
rect 1162 405 1165 413
rect 1179 412 1182 421
rect 1200 424 1203 429
rect 1233 424 1236 429
rect 1200 421 1236 424
rect 1256 424 1259 429
rect 1289 424 1292 429
rect 1256 421 1292 424
rect 1310 424 1313 429
rect 1343 424 1346 429
rect 1310 421 1346 424
rect 1186 412 1189 421
rect 1200 416 1207 417
rect 1200 414 1204 416
rect 1221 412 1225 415
rect 1179 409 1189 412
rect 1162 403 1167 405
rect 1133 395 1136 403
rect 1162 402 1163 403
rect 1179 396 1182 409
rect 1221 408 1224 412
rect 1233 409 1236 421
rect 1289 420 1292 421
rect 1257 413 1260 416
rect 1233 406 1252 409
rect 1233 396 1236 406
rect 1281 410 1284 412
rect 1269 402 1272 408
rect 1283 406 1284 410
rect 1281 405 1284 406
rect 1246 399 1272 402
rect 1289 396 1292 416
rect 1313 412 1314 415
rect 1332 416 1338 417
rect 1332 414 1335 416
rect 1313 403 1316 412
rect 1343 411 1346 421
rect 1315 399 1316 403
rect 1343 396 1346 407
rect 1027 386 1030 392
rect 1099 386 1102 391
rect 1145 386 1148 392
rect 1199 386 1202 392
rect 1255 386 1258 392
rect 1309 386 1312 392
rect 1003 383 1348 386
rect 762 372 964 375
rect 306 371 964 372
rect 306 370 694 371
rect 2 369 229 370
rect 242 369 694 370
rect 2 368 694 369
rect 2 366 367 368
rect 2 362 38 366
rect 42 362 52 366
rect 56 362 66 366
rect 70 363 149 366
rect 70 362 133 363
rect 2 251 6 362
rect 22 361 37 362
rect 36 342 40 349
rect 36 341 41 342
rect 36 337 37 341
rect 44 341 48 362
rect 51 356 64 357
rect 51 352 54 356
rect 58 352 60 356
rect 51 351 64 352
rect 51 344 57 351
rect 67 345 71 362
rect 137 362 149 363
rect 153 363 233 366
rect 153 362 217 363
rect 114 351 126 357
rect 133 356 137 359
rect 221 362 233 363
rect 237 362 270 366
rect 274 362 284 366
rect 288 362 298 366
rect 302 364 367 366
rect 371 364 381 368
rect 385 364 395 368
rect 399 365 478 368
rect 399 364 462 365
rect 302 362 337 364
rect 147 353 169 357
rect 173 353 174 357
rect 198 356 210 357
rect 147 352 151 353
rect 133 351 137 352
rect 114 348 119 351
rect 114 347 115 348
rect 44 337 47 341
rect 51 337 52 341
rect 56 337 57 341
rect 61 337 62 341
rect 67 340 71 341
rect 106 344 115 347
rect 140 348 151 352
rect 198 352 203 356
rect 207 352 210 356
rect 198 351 210 352
rect 217 356 221 359
rect 231 353 253 357
rect 257 353 258 357
rect 231 352 235 353
rect 217 351 221 352
rect 140 344 144 348
rect 158 345 159 349
rect 163 345 174 349
rect 36 336 41 337
rect 36 328 40 336
rect 56 332 62 337
rect 43 328 44 332
rect 48 328 62 332
rect 68 330 72 333
rect 106 330 109 344
rect 114 343 119 344
rect 123 342 144 344
rect 36 319 40 324
rect 36 318 41 319
rect 36 314 37 318
rect 41 314 48 317
rect 36 311 48 314
rect 52 315 56 328
rect 115 338 123 339
rect 127 340 144 342
rect 115 335 127 338
rect 68 324 72 326
rect 59 320 63 324
rect 67 320 72 324
rect 59 319 72 320
rect 115 323 119 335
rect 140 333 144 340
rect 148 338 149 342
rect 153 341 154 342
rect 153 338 165 341
rect 148 337 165 338
rect 161 334 165 337
rect 161 333 166 334
rect 129 327 135 332
rect 140 329 152 333
rect 156 329 157 333
rect 161 329 162 333
rect 129 325 131 327
rect 122 323 131 325
rect 161 328 166 329
rect 170 329 174 345
rect 198 348 203 351
rect 198 344 199 348
rect 224 348 235 352
rect 224 344 228 348
rect 242 345 243 349
rect 247 346 258 349
rect 247 345 261 346
rect 198 343 203 344
rect 207 342 228 344
rect 254 343 261 345
rect 199 338 207 339
rect 211 340 228 342
rect 199 335 211 338
rect 161 324 165 328
rect 122 319 135 323
rect 141 320 165 324
rect 170 325 172 329
rect 115 318 119 319
rect 141 318 145 320
rect 52 311 66 315
rect 70 311 71 315
rect 128 311 129 315
rect 133 311 134 315
rect 170 316 174 325
rect 199 323 203 335
rect 224 333 228 340
rect 232 338 233 342
rect 237 341 238 342
rect 237 338 249 341
rect 232 337 249 338
rect 245 334 249 337
rect 245 333 250 334
rect 213 327 219 332
rect 224 329 236 333
rect 240 329 241 333
rect 245 329 246 333
rect 213 325 215 327
rect 206 323 215 325
rect 245 328 250 329
rect 245 324 249 328
rect 206 319 219 323
rect 225 320 249 324
rect 199 318 203 319
rect 225 318 229 320
rect 141 313 145 314
rect 150 312 151 316
rect 155 312 174 316
rect 128 306 134 311
rect 212 311 213 315
rect 217 311 218 315
rect 254 316 258 343
rect 268 342 272 349
rect 268 341 273 342
rect 268 337 269 341
rect 276 341 280 362
rect 283 356 296 357
rect 283 352 286 356
rect 290 352 292 356
rect 283 351 296 352
rect 283 344 289 351
rect 299 345 303 362
rect 311 343 322 346
rect 276 337 279 341
rect 283 337 284 341
rect 288 337 289 341
rect 293 337 294 341
rect 299 340 303 341
rect 268 336 273 337
rect 268 328 272 336
rect 288 332 294 337
rect 275 328 276 332
rect 280 328 294 332
rect 300 331 304 333
rect 225 313 229 314
rect 234 312 235 316
rect 239 312 258 316
rect 262 325 272 328
rect 262 313 265 325
rect 212 306 218 311
rect 268 319 272 325
rect 268 318 273 319
rect 268 314 269 318
rect 273 314 280 317
rect 268 311 280 314
rect 284 315 288 328
rect 300 324 304 327
rect 291 320 295 324
rect 299 320 304 324
rect 291 319 304 320
rect 284 311 298 315
rect 302 311 303 315
rect 35 302 38 306
rect 42 302 48 306
rect 52 302 116 306
rect 120 302 169 306
rect 173 302 200 306
rect 204 302 253 306
rect 257 302 270 306
rect 274 302 280 306
rect 284 305 308 306
rect 284 302 302 305
rect 21 299 302 302
rect 21 298 308 299
rect 125 296 169 298
rect 125 292 131 296
rect 135 292 159 296
rect 163 292 169 296
rect 129 284 135 292
rect 129 280 130 284
rect 134 280 135 284
rect 140 284 144 285
rect 149 284 155 292
rect 149 280 150 284
rect 154 280 155 284
rect 160 284 165 287
rect 164 280 165 284
rect 140 277 144 280
rect 160 279 165 280
rect 140 273 157 277
rect 129 261 133 271
rect 137 266 142 270
rect 153 269 157 273
rect 137 258 143 262
rect 147 258 150 262
rect 1 231 6 251
rect 137 252 141 258
rect 153 254 157 265
rect 124 249 141 252
rect 145 250 157 254
rect 161 275 322 279
rect 145 246 149 250
rect 161 249 165 275
rect 331 253 335 362
rect 365 344 369 351
rect 365 343 370 344
rect 365 339 366 343
rect 373 343 377 364
rect 380 358 393 359
rect 380 354 383 358
rect 387 354 389 358
rect 380 353 393 354
rect 380 346 386 353
rect 396 347 400 364
rect 466 364 478 365
rect 482 365 562 368
rect 482 364 546 365
rect 443 353 455 359
rect 462 358 466 361
rect 550 364 562 365
rect 566 364 599 368
rect 603 364 613 368
rect 617 364 627 368
rect 631 367 694 368
rect 698 367 708 371
rect 712 367 722 371
rect 726 368 805 371
rect 726 367 789 368
rect 631 364 667 367
rect 476 355 498 359
rect 502 355 503 359
rect 518 358 539 359
rect 476 354 480 355
rect 462 353 466 354
rect 443 350 448 353
rect 373 339 376 343
rect 380 339 381 343
rect 385 339 386 343
rect 390 339 391 343
rect 396 342 400 343
rect 443 349 444 350
rect 365 338 370 339
rect 365 330 369 338
rect 385 334 391 339
rect 372 330 373 334
rect 377 330 391 334
rect 397 332 401 335
rect 365 321 369 326
rect 365 320 370 321
rect 365 316 366 320
rect 370 316 377 319
rect 365 313 377 316
rect 381 317 385 330
rect 397 326 401 328
rect 388 322 392 326
rect 396 322 401 326
rect 388 321 401 322
rect 381 313 395 317
rect 399 313 400 317
rect 418 317 422 345
rect 435 346 444 349
rect 469 350 480 354
rect 518 354 532 358
rect 536 354 539 358
rect 518 353 539 354
rect 546 358 550 361
rect 560 355 582 359
rect 586 355 587 359
rect 560 354 564 355
rect 546 353 550 354
rect 469 346 473 350
rect 487 347 488 351
rect 492 347 503 351
rect 435 332 438 346
rect 443 345 448 346
rect 452 344 473 346
rect 444 340 452 341
rect 456 342 473 344
rect 444 337 456 340
rect 444 325 448 337
rect 469 335 473 342
rect 477 340 478 344
rect 482 343 483 344
rect 482 340 494 343
rect 477 339 494 340
rect 490 336 494 339
rect 490 335 495 336
rect 458 329 464 334
rect 469 331 481 335
rect 485 331 486 335
rect 490 331 491 335
rect 458 327 460 329
rect 451 325 460 327
rect 490 330 495 331
rect 499 331 503 347
rect 527 350 532 353
rect 527 346 528 350
rect 553 350 564 354
rect 553 346 557 350
rect 571 347 572 351
rect 576 347 589 351
rect 527 345 532 346
rect 536 344 557 346
rect 528 340 536 341
rect 540 342 557 344
rect 528 337 540 340
rect 490 326 494 330
rect 451 321 464 325
rect 470 322 494 326
rect 499 327 501 331
rect 444 320 448 321
rect 470 320 474 322
rect 414 314 422 317
rect 457 313 458 317
rect 462 313 463 317
rect 499 318 503 327
rect 528 325 532 337
rect 553 335 557 342
rect 561 340 562 344
rect 566 343 567 344
rect 566 340 578 343
rect 561 339 578 340
rect 574 336 578 339
rect 574 335 579 336
rect 542 329 548 334
rect 553 331 565 335
rect 569 331 570 335
rect 574 331 575 335
rect 542 327 544 329
rect 535 325 544 327
rect 574 330 579 331
rect 574 326 578 330
rect 535 321 548 325
rect 554 322 578 326
rect 528 320 532 321
rect 554 320 558 322
rect 470 315 474 316
rect 479 314 480 318
rect 484 314 503 318
rect 457 308 463 313
rect 541 313 542 317
rect 546 313 547 317
rect 583 318 587 347
rect 597 344 601 351
rect 597 343 602 344
rect 597 339 598 343
rect 605 343 609 364
rect 612 358 625 359
rect 612 354 615 358
rect 619 354 621 358
rect 612 353 625 354
rect 612 346 618 353
rect 628 347 632 364
rect 605 339 608 343
rect 612 339 613 343
rect 617 339 618 343
rect 622 339 623 343
rect 628 342 632 343
rect 597 338 602 339
rect 597 330 601 338
rect 617 334 623 339
rect 604 330 605 334
rect 609 330 623 334
rect 629 333 633 335
rect 554 315 558 316
rect 563 314 564 318
rect 568 314 587 318
rect 591 327 601 330
rect 591 315 594 327
rect 541 308 547 313
rect 597 321 601 327
rect 597 320 602 321
rect 597 316 598 320
rect 602 316 609 319
rect 597 313 609 316
rect 613 317 617 330
rect 629 326 633 329
rect 620 322 624 326
rect 628 322 633 326
rect 620 321 633 322
rect 613 313 627 317
rect 631 313 632 317
rect 364 304 367 308
rect 371 304 377 308
rect 381 304 445 308
rect 449 304 498 308
rect 502 304 529 308
rect 533 304 582 308
rect 586 304 599 308
rect 603 304 609 308
rect 613 307 637 308
rect 613 304 629 307
rect 364 303 629 304
rect 349 301 629 303
rect 635 301 637 307
rect 349 300 637 301
rect 349 299 365 300
rect 454 298 498 300
rect 454 294 460 298
rect 464 294 488 298
rect 492 294 498 298
rect 458 286 464 294
rect 458 282 459 286
rect 463 282 464 286
rect 469 286 473 287
rect 478 286 484 294
rect 478 282 479 286
rect 483 282 484 286
rect 489 286 494 289
rect 584 287 655 290
rect 493 282 494 286
rect 469 279 473 282
rect 489 281 494 282
rect 351 275 419 279
rect 469 275 486 279
rect 458 263 462 273
rect 466 268 471 272
rect 482 271 486 275
rect 466 260 472 264
rect 476 260 479 264
rect 160 248 165 249
rect 129 242 130 246
rect 134 242 149 246
rect 152 244 160 246
rect 164 244 165 248
rect 152 242 165 244
rect 147 236 148 239
rect 125 235 148 236
rect 152 236 153 239
rect 152 235 159 236
rect 125 232 159 235
rect 163 232 169 236
rect 125 231 169 232
rect 330 233 335 253
rect 466 254 470 260
rect 482 256 486 267
rect 453 251 470 254
rect 474 252 486 256
rect 490 275 494 281
rect 490 272 641 275
rect 645 272 646 275
rect 474 248 478 252
rect 490 251 494 272
rect 489 250 494 251
rect 458 244 459 248
rect 463 244 478 248
rect 481 246 489 248
rect 493 246 494 250
rect 481 244 494 246
rect 476 238 477 241
rect 454 237 477 238
rect 481 238 482 241
rect 481 237 488 238
rect 454 234 488 237
rect 492 234 498 238
rect 454 233 498 234
rect 1 228 169 231
rect 1 227 129 228
rect 307 227 322 231
rect 126 224 129 227
rect 330 230 498 233
rect 330 229 456 230
rect 453 226 456 229
rect 1 220 307 224
rect 1 216 37 220
rect 41 216 51 220
rect 55 216 65 220
rect 69 217 148 220
rect 69 216 132 217
rect 1 105 5 216
rect 35 196 39 203
rect 35 195 40 196
rect 35 191 36 195
rect 43 195 47 216
rect 50 210 63 211
rect 50 206 53 210
rect 57 206 59 210
rect 50 205 63 206
rect 50 198 56 205
rect 66 199 70 216
rect 136 216 148 217
rect 152 217 232 220
rect 152 216 216 217
rect 113 205 125 211
rect 132 210 136 213
rect 220 216 232 217
rect 236 216 269 220
rect 273 216 283 220
rect 287 216 297 220
rect 301 216 307 220
rect 330 222 636 226
rect 651 225 654 287
rect 658 256 662 364
rect 692 347 696 354
rect 692 346 697 347
rect 692 342 693 346
rect 700 346 704 367
rect 707 361 720 362
rect 707 357 710 361
rect 714 357 716 361
rect 707 356 720 357
rect 707 349 713 356
rect 723 350 727 367
rect 793 367 805 368
rect 809 368 889 371
rect 809 367 873 368
rect 770 356 782 362
rect 789 361 793 364
rect 877 367 889 368
rect 893 367 926 371
rect 930 367 940 371
rect 944 367 954 371
rect 958 367 964 371
rect 803 358 825 362
rect 829 358 830 362
rect 843 361 866 362
rect 803 357 807 358
rect 843 357 859 361
rect 863 357 866 361
rect 789 356 793 357
rect 770 353 775 356
rect 770 352 771 353
rect 700 342 703 346
rect 707 342 708 346
rect 712 342 713 346
rect 717 342 718 346
rect 723 345 727 346
rect 692 341 697 342
rect 692 333 696 341
rect 712 337 718 342
rect 699 333 700 337
rect 704 333 718 337
rect 724 335 728 338
rect 692 324 696 329
rect 692 323 697 324
rect 692 319 693 323
rect 697 319 704 322
rect 692 316 704 319
rect 708 320 712 333
rect 724 329 728 331
rect 715 325 719 329
rect 723 325 728 329
rect 715 324 728 325
rect 708 316 722 320
rect 726 316 727 320
rect 751 318 755 347
rect 762 349 771 352
rect 796 353 807 357
rect 796 349 800 353
rect 814 350 815 354
rect 819 350 830 354
rect 762 335 765 349
rect 770 348 775 349
rect 779 347 800 349
rect 771 343 779 344
rect 783 345 800 347
rect 771 340 783 343
rect 771 328 775 340
rect 796 338 800 345
rect 804 343 805 347
rect 809 346 810 347
rect 809 343 821 346
rect 804 342 821 343
rect 817 339 821 342
rect 817 338 822 339
rect 785 332 791 337
rect 796 334 808 338
rect 812 334 813 338
rect 817 334 818 338
rect 785 330 787 332
rect 778 328 787 330
rect 817 333 822 334
rect 826 334 830 350
rect 817 329 821 333
rect 778 324 791 328
rect 797 325 821 329
rect 826 330 828 334
rect 771 323 775 324
rect 797 323 801 325
rect 751 314 752 318
rect 784 316 785 320
rect 789 316 790 320
rect 826 321 830 330
rect 797 318 801 319
rect 806 317 807 321
rect 811 317 830 321
rect 837 318 840 349
rect 784 311 790 316
rect 844 311 848 357
rect 854 356 866 357
rect 873 361 877 364
rect 887 358 909 362
rect 913 358 914 362
rect 887 357 891 358
rect 873 356 877 357
rect 854 353 859 356
rect 854 349 855 353
rect 880 353 891 357
rect 880 349 884 353
rect 898 350 899 354
rect 903 350 914 354
rect 854 348 859 349
rect 863 347 884 349
rect 855 343 863 344
rect 867 345 884 347
rect 855 340 867 343
rect 855 328 859 340
rect 880 338 884 345
rect 888 343 889 347
rect 893 346 894 347
rect 893 343 905 346
rect 888 342 905 343
rect 901 339 905 342
rect 901 338 906 339
rect 869 332 875 337
rect 880 334 892 338
rect 896 334 897 338
rect 901 334 902 338
rect 869 330 871 332
rect 862 328 871 330
rect 901 333 906 334
rect 901 329 905 333
rect 862 324 875 328
rect 881 325 905 329
rect 855 323 859 324
rect 881 323 885 325
rect 868 316 869 320
rect 873 316 874 320
rect 910 321 914 350
rect 924 347 928 354
rect 924 346 929 347
rect 924 342 925 346
rect 932 346 936 367
rect 939 361 952 362
rect 939 357 942 361
rect 946 357 948 361
rect 939 356 952 357
rect 939 349 945 356
rect 955 350 959 367
rect 932 342 935 346
rect 939 342 940 346
rect 944 342 945 346
rect 949 342 950 346
rect 955 345 959 346
rect 924 341 929 342
rect 924 333 928 341
rect 944 337 950 342
rect 931 333 932 337
rect 936 333 950 337
rect 956 336 960 338
rect 881 318 885 319
rect 890 317 891 321
rect 895 317 914 321
rect 918 330 928 333
rect 918 318 921 330
rect 868 311 874 316
rect 924 324 928 330
rect 924 323 929 324
rect 924 319 925 323
rect 929 319 936 322
rect 924 316 936 319
rect 940 320 944 333
rect 956 329 960 332
rect 1003 330 1007 383
rect 1171 380 1176 383
rect 1277 380 1281 383
rect 1103 377 1352 380
rect 1103 372 1106 377
rect 1149 371 1152 377
rect 1203 371 1206 377
rect 1259 371 1262 377
rect 1313 371 1316 377
rect 1137 360 1140 368
rect 1137 356 1138 360
rect 947 325 951 329
rect 955 325 960 329
rect 947 324 960 325
rect 971 326 1007 330
rect 940 316 954 320
rect 958 316 959 320
rect 691 310 694 311
rect 689 307 694 310
rect 698 307 704 311
rect 708 307 772 311
rect 776 307 825 311
rect 829 307 856 311
rect 860 307 909 311
rect 913 307 926 311
rect 930 307 936 311
rect 940 307 964 311
rect 971 307 975 326
rect 689 305 975 307
rect 676 303 975 305
rect 676 302 693 303
rect 676 301 692 302
rect 781 301 825 303
rect 781 297 787 301
rect 791 297 815 301
rect 819 297 825 301
rect 785 289 791 297
rect 785 285 786 289
rect 790 285 791 289
rect 796 289 800 290
rect 805 289 811 297
rect 805 285 806 289
rect 810 285 811 289
rect 816 289 821 292
rect 820 285 821 289
rect 677 272 744 275
rect 748 272 749 275
rect 657 236 662 256
rect 754 244 758 284
rect 796 282 800 285
rect 816 284 821 285
rect 796 278 813 282
rect 766 250 769 277
rect 785 266 789 276
rect 793 271 798 275
rect 809 274 813 278
rect 793 263 799 267
rect 803 263 806 267
rect 793 257 797 263
rect 809 259 813 270
rect 780 254 797 257
rect 801 255 813 259
rect 817 280 821 284
rect 817 277 829 280
rect 801 251 805 255
rect 817 254 821 277
rect 837 256 840 271
rect 816 253 821 254
rect 785 247 786 251
rect 790 247 805 251
rect 808 249 816 251
rect 820 249 821 253
rect 808 247 821 249
rect 803 241 804 244
rect 754 239 758 240
rect 781 240 804 241
rect 808 241 809 244
rect 836 243 841 256
rect 808 240 815 241
rect 781 237 815 240
rect 819 237 825 241
rect 781 236 825 237
rect 987 241 990 326
rect 1086 322 1090 350
rect 1120 347 1123 350
rect 1137 334 1140 356
rect 1183 354 1186 367
rect 1183 351 1193 354
rect 1225 351 1228 355
rect 1237 357 1240 367
rect 1237 354 1256 357
rect 1285 357 1288 358
rect 1152 347 1154 350
rect 1174 347 1175 350
rect 1183 342 1186 351
rect 1150 339 1186 342
rect 1150 334 1153 339
rect 1183 334 1186 339
rect 1190 342 1193 351
rect 1204 347 1208 349
rect 1225 348 1229 351
rect 1204 346 1211 347
rect 1237 342 1240 354
rect 1287 353 1288 357
rect 1285 351 1288 353
rect 1261 347 1264 350
rect 1293 347 1296 367
rect 1319 360 1320 364
rect 1317 351 1320 360
rect 1347 356 1350 367
rect 1317 348 1318 351
rect 1336 347 1339 349
rect 1336 346 1342 347
rect 1293 342 1296 343
rect 1347 342 1350 352
rect 1204 339 1240 342
rect 1204 334 1207 339
rect 1237 334 1240 339
rect 1260 339 1296 342
rect 1260 334 1263 339
rect 1293 334 1296 339
rect 1314 339 1350 342
rect 1314 334 1317 339
rect 1347 334 1350 339
rect 1089 320 1090 322
rect 1103 311 1106 330
rect 1166 311 1169 330
rect 1176 311 1179 316
rect 1220 311 1223 330
rect 1230 311 1233 316
rect 1276 311 1279 330
rect 1286 311 1289 316
rect 1330 311 1333 330
rect 1340 311 1343 316
rect 1361 311 1366 452
rect 1496 356 1500 475
rect 1631 473 1655 475
rect 1631 472 1672 473
rect 1631 468 1651 472
rect 1655 469 1672 472
rect 1676 469 1677 473
rect 1684 470 1686 474
rect 1690 470 1698 474
rect 1693 469 1698 470
rect 1560 371 1563 463
rect 1631 458 1655 468
rect 1631 454 1651 458
rect 1631 450 1655 454
rect 1660 462 1661 466
rect 1665 462 1666 466
rect 1697 465 1698 469
rect 1660 460 1666 462
rect 1660 456 1661 460
rect 1665 459 1666 460
rect 1676 463 1689 464
rect 1680 459 1689 463
rect 1693 461 1698 465
rect 1702 472 1706 473
rect 1665 456 1673 459
rect 1676 458 1689 459
rect 1702 458 1706 468
rect 1660 453 1673 456
rect 1685 454 1706 458
rect 1711 454 1719 478
rect 1676 453 1680 454
rect 1631 449 1676 450
rect 1631 446 1680 449
rect 1685 450 1689 454
rect 1715 450 1719 454
rect 1567 443 1575 446
rect 1567 439 1571 443
rect 1567 433 1575 439
rect 1580 444 1593 445
rect 1580 440 1583 444
rect 1587 441 1593 444
rect 1597 444 1618 445
rect 1597 441 1606 444
rect 1587 440 1588 441
rect 1605 440 1606 441
rect 1610 441 1618 444
rect 1631 444 1655 446
rect 1685 445 1689 446
rect 1631 443 1651 444
rect 1610 440 1611 441
rect 1580 433 1586 440
rect 1635 440 1651 443
rect 1700 443 1706 450
rect 1675 442 1676 443
rect 1635 439 1655 440
rect 1597 437 1601 438
rect 1631 437 1655 439
rect 1668 439 1676 442
rect 1680 442 1681 443
rect 1698 442 1699 443
rect 1680 439 1699 442
rect 1703 439 1706 443
rect 1668 438 1706 439
rect 1711 444 1719 450
rect 1715 440 1719 444
rect 1567 429 1571 433
rect 1597 429 1601 433
rect 1606 434 1655 437
rect 1610 433 1655 434
rect 1689 435 1692 438
rect 1606 429 1610 430
rect 1567 365 1575 429
rect 1580 425 1601 429
rect 1613 427 1626 430
rect 1580 415 1584 425
rect 1597 424 1610 425
rect 1613 424 1621 427
rect 1580 410 1584 411
rect 1588 418 1593 422
rect 1597 420 1606 424
rect 1597 419 1610 420
rect 1620 423 1621 424
rect 1625 423 1626 427
rect 1620 421 1626 423
rect 1588 414 1589 418
rect 1620 417 1621 421
rect 1625 417 1626 421
rect 1631 429 1655 433
rect 1635 425 1655 429
rect 1689 432 1704 435
rect 1676 428 1680 429
rect 1631 415 1655 425
rect 1588 413 1593 414
rect 1588 409 1595 413
rect 1599 409 1602 413
rect 1609 410 1610 414
rect 1614 411 1631 414
rect 1635 411 1655 415
rect 1614 410 1655 411
rect 1631 407 1655 410
rect 1631 403 1651 407
rect 1585 396 1621 399
rect 1631 391 1655 403
rect 1660 427 1664 428
rect 1660 405 1664 423
rect 1668 424 1705 428
rect 1668 417 1672 424
rect 1683 419 1684 420
rect 1668 412 1672 413
rect 1676 416 1684 419
rect 1688 419 1689 420
rect 1688 416 1697 419
rect 1676 415 1697 416
rect 1676 408 1680 415
rect 1675 407 1680 408
rect 1660 401 1669 405
rect 1679 403 1680 407
rect 1675 402 1680 403
rect 1684 410 1688 411
rect 1665 398 1669 401
rect 1684 398 1688 406
rect 1665 394 1688 398
rect 1693 399 1697 415
rect 1701 409 1705 424
rect 1701 404 1705 405
rect 1711 427 1719 440
rect 1715 423 1719 427
rect 1693 395 1699 399
rect 1703 395 1704 399
rect 1631 387 1654 391
rect 1658 387 1661 391
rect 1665 387 1666 391
rect 1599 372 1616 375
rect 1613 367 1616 372
rect 1612 366 1626 367
rect 1567 361 1571 365
rect 1587 362 1588 366
rect 1592 362 1608 366
rect 1612 362 1613 366
rect 1617 362 1626 366
rect 1497 334 1505 356
rect 1511 351 1515 352
rect 1511 336 1515 347
rect 1518 344 1521 357
rect 1567 356 1575 361
rect 1561 353 1575 356
rect 1561 352 1584 353
rect 1530 348 1540 352
rect 1549 351 1580 352
rect 1553 350 1580 351
rect 1553 347 1561 350
rect 1549 346 1561 347
rect 1565 348 1580 350
rect 1565 347 1584 348
rect 1588 352 1594 359
rect 1604 358 1608 362
rect 1604 354 1607 358
rect 1611 354 1613 358
rect 1620 355 1626 362
rect 1588 350 1601 352
rect 1565 346 1575 347
rect 1588 346 1592 350
rect 1596 346 1601 350
rect 1518 340 1531 344
rect 1527 338 1531 340
rect 1535 339 1539 344
rect 1497 333 1508 334
rect 1497 329 1504 333
rect 1511 332 1523 336
rect 1497 328 1508 329
rect 1497 322 1505 328
rect 1497 318 1501 322
rect 1497 312 1505 318
rect 1511 321 1515 329
rect 1519 328 1523 332
rect 1542 337 1549 341
rect 1553 337 1554 341
rect 1527 331 1531 334
rect 1542 328 1546 337
rect 1561 332 1575 346
rect 1609 341 1613 354
rect 1631 348 1655 387
rect 1673 381 1677 394
rect 1685 385 1690 389
rect 1694 385 1698 389
rect 1711 388 1719 423
rect 1685 383 1698 385
rect 1660 377 1666 380
rect 1673 377 1675 381
rect 1679 377 1682 381
rect 1660 373 1661 377
rect 1665 373 1666 377
rect 1678 373 1682 377
rect 1692 376 1698 383
rect 1702 387 1719 388
rect 1706 383 1719 387
rect 1702 382 1719 383
rect 1711 374 1719 382
rect 1660 369 1669 373
rect 1673 369 1674 373
rect 1678 369 1694 373
rect 1698 369 1699 373
rect 1715 370 1719 374
rect 1660 368 1674 369
rect 1664 354 1703 357
rect 1707 354 1708 357
rect 1620 344 1621 348
rect 1625 344 1628 348
rect 1632 344 1655 348
rect 1582 336 1583 340
rect 1587 336 1593 340
rect 1519 324 1534 328
rect 1538 324 1546 328
rect 1549 331 1575 332
rect 1553 327 1575 331
rect 1549 326 1575 327
rect 1561 322 1575 326
rect 1511 317 1513 321
rect 1517 320 1518 321
rect 1548 320 1549 321
rect 1517 317 1549 320
rect 1553 317 1556 321
rect 1511 316 1556 317
rect 1565 318 1575 322
rect 1101 310 1366 311
rect 1000 307 1408 310
rect 1016 288 1019 307
rect 1099 288 1102 307
rect 1112 299 1142 302
rect 1061 273 1065 284
rect 1044 269 1047 272
rect 1061 263 1064 273
rect 1116 268 1119 271
rect 1061 259 1062 263
rect 1133 262 1136 284
rect 1139 272 1142 299
rect 1162 288 1165 307
rect 1172 302 1175 307
rect 1216 288 1219 307
rect 1226 302 1229 307
rect 1272 288 1275 307
rect 1282 302 1285 307
rect 1326 288 1329 307
rect 1336 302 1339 307
rect 1146 279 1149 284
rect 1179 279 1182 284
rect 1146 276 1182 279
rect 1139 269 1144 272
rect 1148 268 1150 271
rect 1170 268 1171 271
rect 1179 267 1182 276
rect 1200 279 1203 284
rect 1233 279 1236 284
rect 1200 276 1236 279
rect 1256 279 1259 284
rect 1289 279 1292 284
rect 1256 276 1292 279
rect 1310 279 1313 284
rect 1343 279 1346 284
rect 1310 276 1346 279
rect 1186 267 1189 276
rect 1200 271 1207 272
rect 1200 269 1204 271
rect 1221 267 1225 270
rect 1179 264 1189 267
rect 1061 251 1064 259
rect 1133 258 1134 262
rect 1133 250 1136 258
rect 1179 251 1182 264
rect 1221 263 1224 267
rect 1233 264 1236 276
rect 1289 275 1292 276
rect 1257 268 1260 271
rect 1233 261 1252 264
rect 1233 251 1236 261
rect 1281 265 1284 267
rect 1269 257 1272 263
rect 1283 261 1284 265
rect 1281 260 1284 261
rect 1246 254 1272 257
rect 1289 251 1292 271
rect 1313 267 1314 270
rect 1332 271 1338 272
rect 1332 269 1335 271
rect 1313 258 1316 267
rect 1343 266 1346 276
rect 1315 254 1316 258
rect 1343 251 1346 262
rect 1027 241 1030 247
rect 1099 241 1102 246
rect 1145 241 1148 247
rect 1199 241 1202 247
rect 1255 241 1258 247
rect 1309 241 1312 247
rect 959 237 981 240
rect 657 233 825 236
rect 657 232 781 233
rect 786 229 789 233
rect 330 218 366 222
rect 370 218 380 222
rect 384 218 394 222
rect 398 219 477 222
rect 398 218 461 219
rect 146 207 168 211
rect 172 207 173 211
rect 197 210 209 211
rect 185 207 202 210
rect 146 206 150 207
rect 132 205 136 206
rect 113 202 118 205
rect 113 201 114 202
rect 43 191 46 195
rect 50 191 51 195
rect 55 191 56 195
rect 60 191 61 195
rect 66 194 70 195
rect 105 198 114 201
rect 139 202 150 206
rect 139 198 143 202
rect 157 199 158 203
rect 162 199 173 203
rect 35 190 40 191
rect 35 182 39 190
rect 55 186 61 191
rect 42 182 43 186
rect 47 182 61 186
rect 67 184 71 187
rect 105 184 108 198
rect 113 197 118 198
rect 122 196 143 198
rect 35 173 39 178
rect 35 172 40 173
rect 35 168 36 172
rect 40 168 47 171
rect 35 165 47 168
rect 51 169 55 182
rect 114 192 122 193
rect 126 194 143 196
rect 114 189 126 192
rect 67 178 71 180
rect 58 174 62 178
rect 66 174 71 178
rect 58 173 71 174
rect 114 177 118 189
rect 139 187 143 194
rect 147 192 148 196
rect 152 195 153 196
rect 152 192 164 195
rect 147 191 164 192
rect 160 188 164 191
rect 160 187 165 188
rect 128 181 134 186
rect 139 183 151 187
rect 155 183 156 187
rect 160 183 161 187
rect 128 179 130 181
rect 121 177 130 179
rect 160 182 165 183
rect 169 183 173 199
rect 160 178 164 182
rect 121 173 134 177
rect 140 174 164 178
rect 169 179 171 183
rect 114 172 118 173
rect 140 172 144 174
rect 51 165 65 169
rect 69 165 70 169
rect 127 165 128 169
rect 132 165 133 169
rect 169 170 173 179
rect 140 167 144 168
rect 149 166 150 170
rect 154 166 173 170
rect 185 167 188 207
rect 197 206 202 207
rect 206 206 209 210
rect 197 205 209 206
rect 216 210 220 213
rect 230 207 252 211
rect 256 207 257 211
rect 230 206 234 207
rect 216 205 220 206
rect 197 202 202 205
rect 197 198 198 202
rect 223 202 234 206
rect 223 198 227 202
rect 241 199 242 203
rect 246 199 257 203
rect 197 197 202 198
rect 206 196 227 198
rect 198 192 206 193
rect 210 194 227 196
rect 198 189 210 192
rect 198 177 202 189
rect 223 187 227 194
rect 231 192 232 196
rect 236 195 237 196
rect 236 192 248 195
rect 231 191 248 192
rect 244 188 248 191
rect 253 191 257 199
rect 267 196 271 203
rect 267 195 272 196
rect 267 191 268 195
rect 275 195 279 216
rect 282 210 295 211
rect 282 206 285 210
rect 289 206 291 210
rect 282 205 295 206
rect 282 198 288 205
rect 298 199 302 216
rect 312 198 327 201
rect 275 191 278 195
rect 282 191 283 195
rect 287 191 288 195
rect 292 191 293 195
rect 298 194 302 195
rect 244 187 249 188
rect 212 181 218 186
rect 223 183 235 187
rect 239 183 240 187
rect 244 183 245 187
rect 212 179 214 181
rect 205 177 214 179
rect 244 182 249 183
rect 253 187 260 191
rect 267 190 272 191
rect 244 178 248 182
rect 205 173 218 177
rect 224 174 248 178
rect 198 172 202 173
rect 224 172 228 174
rect 127 160 133 165
rect 211 165 212 169
rect 216 165 217 169
rect 253 170 257 187
rect 267 182 271 190
rect 287 186 293 191
rect 274 182 275 186
rect 279 182 293 186
rect 299 185 303 187
rect 224 167 228 168
rect 233 166 234 170
rect 238 166 257 170
rect 261 179 271 182
rect 261 167 264 179
rect 211 160 217 165
rect 267 173 271 179
rect 267 172 272 173
rect 267 168 268 172
rect 272 168 279 171
rect 267 165 279 168
rect 283 169 287 182
rect 299 178 303 181
rect 290 174 294 178
rect 298 174 303 178
rect 290 173 303 174
rect 283 165 297 169
rect 301 165 302 169
rect 34 156 37 160
rect 41 156 47 160
rect 51 156 115 160
rect 119 156 168 160
rect 172 156 199 160
rect 203 156 252 160
rect 256 156 269 160
rect 273 156 279 160
rect 283 156 302 160
rect 34 153 302 156
rect 34 152 307 153
rect 124 150 168 152
rect 124 146 130 150
rect 134 146 158 150
rect 162 146 168 150
rect 324 148 327 198
rect 128 138 134 146
rect 128 134 129 138
rect 133 134 134 138
rect 139 138 143 139
rect 148 138 154 146
rect 255 143 296 146
rect 325 144 327 148
rect 148 134 149 138
rect 153 134 154 138
rect 159 138 164 141
rect 163 134 164 138
rect 139 131 143 134
rect 159 133 164 134
rect 139 127 156 131
rect 128 115 132 125
rect 136 120 141 124
rect 152 123 156 127
rect 136 112 142 116
rect 146 112 149 116
rect 0 87 5 105
rect 136 106 140 112
rect 152 108 156 119
rect 123 103 140 106
rect 144 104 156 108
rect 160 122 164 133
rect 252 125 275 128
rect 280 125 281 128
rect 160 119 187 122
rect 144 100 148 104
rect 160 103 164 119
rect 159 102 164 103
rect 128 96 129 100
rect 133 96 148 100
rect 151 98 159 100
rect 163 98 164 102
rect 151 96 164 98
rect 181 109 187 119
rect 146 90 147 93
rect -37 85 5 87
rect 124 89 147 90
rect 151 90 152 93
rect 151 89 158 90
rect 124 86 158 89
rect 162 86 168 90
rect 124 85 168 86
rect -37 82 168 85
rect -37 81 124 82
rect -37 80 4 81
rect -37 76 -31 80
rect -36 -134 -31 76
rect 181 13 188 109
rect 293 42 296 143
rect 305 124 321 128
rect 330 107 334 218
rect 364 198 368 205
rect 364 197 369 198
rect 364 193 365 197
rect 372 197 376 218
rect 379 212 392 213
rect 379 208 382 212
rect 386 208 388 212
rect 379 207 392 208
rect 379 200 385 207
rect 395 201 399 218
rect 465 218 477 219
rect 481 219 561 222
rect 481 218 545 219
rect 442 207 454 213
rect 461 212 465 215
rect 549 218 561 219
rect 565 218 598 222
rect 602 218 612 222
rect 616 218 626 222
rect 630 218 636 222
rect 650 222 654 225
rect 657 225 963 229
rect 475 209 497 213
rect 501 209 502 213
rect 526 212 538 213
rect 475 208 479 209
rect 461 207 465 208
rect 442 204 447 207
rect 442 203 443 204
rect 372 193 375 197
rect 379 193 380 197
rect 384 193 385 197
rect 389 193 390 197
rect 395 196 399 197
rect 434 200 443 203
rect 468 204 479 208
rect 526 208 531 212
rect 535 208 538 212
rect 526 207 538 208
rect 545 212 549 215
rect 559 209 581 213
rect 585 209 586 213
rect 559 208 563 209
rect 545 207 549 208
rect 468 200 472 204
rect 486 201 487 205
rect 491 201 502 205
rect 364 192 369 193
rect 364 184 368 192
rect 384 188 390 193
rect 371 184 372 188
rect 376 184 390 188
rect 396 186 400 189
rect 364 175 368 180
rect 364 174 369 175
rect 364 170 365 174
rect 369 170 376 173
rect 364 167 376 170
rect 380 171 384 184
rect 396 180 400 182
rect 387 176 391 180
rect 395 176 400 180
rect 387 175 400 176
rect 380 167 394 171
rect 398 167 399 171
rect 424 169 427 189
rect 434 186 437 200
rect 442 199 447 200
rect 451 198 472 200
rect 443 194 451 195
rect 455 196 472 198
rect 443 191 455 194
rect 443 179 447 191
rect 468 189 472 196
rect 476 194 477 198
rect 481 197 482 198
rect 481 194 493 197
rect 476 193 493 194
rect 489 190 493 193
rect 489 189 494 190
rect 457 183 463 188
rect 468 185 480 189
rect 484 185 485 189
rect 489 185 490 189
rect 457 181 459 183
rect 450 179 459 181
rect 489 184 494 185
rect 498 185 502 201
rect 526 204 531 207
rect 526 200 527 204
rect 552 204 563 208
rect 552 200 556 204
rect 570 201 571 205
rect 575 201 586 205
rect 526 199 531 200
rect 535 198 556 200
rect 527 194 535 195
rect 539 196 556 198
rect 527 191 539 194
rect 489 180 493 184
rect 450 175 463 179
rect 469 176 493 180
rect 498 181 500 185
rect 443 174 447 175
rect 469 174 473 176
rect 456 167 457 171
rect 461 167 462 171
rect 498 172 502 181
rect 527 179 531 191
rect 552 189 556 196
rect 560 194 561 198
rect 565 197 566 198
rect 565 194 577 197
rect 560 193 577 194
rect 573 190 577 193
rect 582 196 586 201
rect 596 198 600 205
rect 596 197 601 198
rect 582 193 589 196
rect 596 193 597 197
rect 604 197 608 218
rect 611 212 624 213
rect 611 208 614 212
rect 618 208 620 212
rect 611 207 624 208
rect 611 200 617 207
rect 627 201 631 218
rect 604 193 607 197
rect 611 193 612 197
rect 616 193 617 197
rect 621 193 622 197
rect 627 196 631 197
rect 573 189 578 190
rect 541 183 547 188
rect 552 185 564 189
rect 568 185 569 189
rect 573 185 574 189
rect 541 181 543 183
rect 534 179 543 181
rect 573 184 578 185
rect 573 180 577 184
rect 534 175 547 179
rect 553 176 577 180
rect 527 174 531 175
rect 553 174 557 176
rect 469 169 473 170
rect 478 168 479 172
rect 483 168 502 172
rect 456 162 462 167
rect 540 167 541 171
rect 545 167 546 171
rect 582 172 586 193
rect 596 192 601 193
rect 596 184 600 192
rect 616 188 622 193
rect 603 184 604 188
rect 608 184 622 188
rect 628 187 632 189
rect 553 169 557 170
rect 562 168 563 172
rect 567 168 586 172
rect 590 181 600 184
rect 590 169 593 181
rect 540 162 546 167
rect 596 175 600 181
rect 596 174 601 175
rect 596 170 597 174
rect 601 170 608 173
rect 596 167 608 170
rect 612 171 616 184
rect 650 186 653 222
rect 628 180 632 183
rect 619 176 623 180
rect 627 176 632 180
rect 619 175 632 176
rect 648 179 653 186
rect 657 221 693 225
rect 697 221 707 225
rect 711 221 721 225
rect 725 222 804 225
rect 725 221 788 222
rect 612 167 626 171
rect 630 167 631 171
rect 363 158 366 162
rect 370 158 376 162
rect 380 158 444 162
rect 448 158 497 162
rect 501 158 528 162
rect 532 158 581 162
rect 585 158 598 162
rect 602 158 608 162
rect 612 158 636 162
rect 344 155 629 158
rect 363 154 629 155
rect 633 154 636 158
rect 453 152 497 154
rect 453 148 459 152
rect 463 148 487 152
rect 491 148 497 152
rect 352 144 373 147
rect 329 87 334 107
rect 369 109 372 144
rect 424 143 427 145
rect 457 140 463 148
rect 424 125 427 139
rect 457 136 458 140
rect 462 136 463 140
rect 468 140 472 141
rect 477 140 483 148
rect 623 143 627 144
rect 648 143 652 179
rect 477 136 478 140
rect 482 136 483 140
rect 488 140 493 143
rect 492 136 493 140
rect 623 140 652 143
rect 623 139 650 140
rect 468 133 472 136
rect 488 135 493 136
rect 468 129 485 133
rect 396 121 424 124
rect 369 106 389 109
rect 386 97 389 106
rect 383 95 389 97
rect 387 93 389 95
rect 396 95 400 121
rect 457 117 461 127
rect 465 122 470 126
rect 481 125 485 129
rect 465 114 471 118
rect 475 114 478 118
rect 465 108 469 114
rect 481 110 485 121
rect 452 105 469 108
rect 473 106 485 110
rect 473 102 477 106
rect 489 105 493 135
rect 520 131 602 136
rect 623 116 627 139
rect 488 104 493 105
rect 457 98 458 102
rect 462 98 477 102
rect 480 100 488 102
rect 492 102 493 104
rect 492 100 497 102
rect 480 98 497 100
rect 475 92 476 95
rect 453 91 476 92
rect 480 92 481 95
rect 480 91 487 92
rect 453 88 487 91
rect 491 88 497 92
rect 453 87 497 88
rect 329 84 497 87
rect 329 83 377 84
rect 395 83 401 84
rect 419 83 453 84
rect 389 77 407 80
rect 442 76 446 83
rect 325 74 369 76
rect 418 74 462 76
rect 505 74 549 76
rect 325 72 549 74
rect 325 68 331 72
rect 335 71 424 72
rect 335 68 369 71
rect 418 68 424 71
rect 428 71 511 72
rect 428 68 462 71
rect 505 68 511 71
rect 515 68 549 72
rect 339 60 345 68
rect 339 56 340 60
rect 344 56 345 60
rect 350 62 354 63
rect 359 62 365 68
rect 400 62 411 65
rect 359 58 360 62
rect 364 58 365 62
rect 329 55 334 56
rect 329 51 330 55
rect 350 55 354 58
rect 329 48 334 51
rect 329 44 330 48
rect 329 43 334 44
rect 337 51 350 53
rect 337 49 354 51
rect 361 51 392 55
rect 329 42 333 43
rect 293 38 333 42
rect 329 25 333 38
rect 337 38 341 49
rect 352 42 357 46
rect 361 42 365 51
rect 344 34 347 38
rect 351 34 358 38
rect 337 30 341 34
rect 337 26 349 30
rect 353 29 358 34
rect 329 24 334 25
rect 329 20 330 24
rect 334 20 341 23
rect 329 17 341 20
rect 345 22 349 26
rect 352 25 368 29
rect 345 18 360 22
rect 364 18 365 22
rect 388 18 392 51
rect 408 52 411 62
rect 432 60 438 68
rect 432 56 433 60
rect 437 56 438 60
rect 443 62 447 63
rect 452 62 458 68
rect 452 58 453 62
rect 457 58 458 62
rect 519 60 525 68
rect 498 59 514 60
rect 422 55 427 56
rect 422 52 423 55
rect 408 51 423 52
rect 443 55 447 58
rect 408 49 427 51
rect 422 48 427 49
rect 422 44 423 48
rect 422 43 427 44
rect 430 51 443 53
rect 430 49 447 51
rect 422 25 426 43
rect 430 38 434 49
rect 454 46 458 55
rect 502 55 514 59
rect 519 56 520 60
rect 524 56 525 60
rect 530 62 534 63
rect 539 62 545 68
rect 539 58 540 62
rect 544 58 545 62
rect 502 54 510 55
rect 509 51 510 54
rect 530 55 534 58
rect 509 48 514 51
rect 445 42 450 46
rect 454 42 465 46
rect 509 44 510 48
rect 509 43 514 44
rect 517 51 530 53
rect 517 49 534 51
rect 437 34 440 38
rect 444 34 451 38
rect 430 30 434 34
rect 430 26 442 30
rect 422 24 427 25
rect 422 20 423 24
rect 427 20 434 23
rect 422 17 434 20
rect 438 22 442 26
rect 446 29 451 34
rect 446 25 461 29
rect 509 25 513 43
rect 517 38 521 49
rect 541 46 545 55
rect 532 42 537 46
rect 541 42 554 46
rect 585 38 589 76
rect 622 78 627 116
rect 657 110 661 221
rect 691 201 695 208
rect 691 200 696 201
rect 691 196 692 200
rect 699 200 703 221
rect 706 215 719 216
rect 706 211 709 215
rect 713 211 715 215
rect 706 210 719 211
rect 706 203 712 210
rect 722 204 726 221
rect 792 221 804 222
rect 808 222 888 225
rect 808 221 872 222
rect 769 210 781 216
rect 788 215 792 218
rect 876 221 888 222
rect 892 221 925 225
rect 929 221 939 225
rect 943 221 953 225
rect 957 221 963 225
rect 802 212 824 216
rect 828 212 829 216
rect 853 215 865 216
rect 802 211 806 212
rect 788 210 792 211
rect 769 207 774 210
rect 769 206 770 207
rect 699 196 702 200
rect 706 196 707 200
rect 711 196 712 200
rect 716 196 717 200
rect 722 199 726 200
rect 761 203 770 206
rect 795 207 806 211
rect 853 211 858 215
rect 862 211 865 215
rect 853 210 865 211
rect 872 215 876 218
rect 886 212 908 216
rect 912 212 913 216
rect 886 211 890 212
rect 872 210 876 211
rect 795 203 799 207
rect 813 204 814 208
rect 818 204 829 208
rect 691 195 696 196
rect 691 187 695 195
rect 711 191 717 196
rect 698 187 699 191
rect 703 187 717 191
rect 723 189 727 192
rect 761 189 764 203
rect 769 202 774 203
rect 778 201 799 203
rect 691 178 695 183
rect 691 177 696 178
rect 691 173 692 177
rect 696 173 703 176
rect 691 170 703 173
rect 707 174 711 187
rect 770 197 778 198
rect 782 199 799 201
rect 770 194 782 197
rect 723 183 727 185
rect 714 179 718 183
rect 722 179 727 183
rect 714 178 727 179
rect 770 182 774 194
rect 795 192 799 199
rect 803 197 804 201
rect 808 200 809 201
rect 808 197 820 200
rect 803 196 820 197
rect 816 193 820 196
rect 816 192 821 193
rect 784 186 790 191
rect 795 188 807 192
rect 811 188 812 192
rect 816 188 817 192
rect 784 184 786 186
rect 770 177 774 178
rect 777 182 786 184
rect 816 187 821 188
rect 825 188 829 204
rect 853 207 858 210
rect 853 203 854 207
rect 879 207 890 211
rect 879 203 883 207
rect 897 204 898 208
rect 902 204 913 208
rect 853 202 858 203
rect 862 201 883 203
rect 854 197 862 198
rect 866 199 883 201
rect 854 194 866 197
rect 816 183 820 187
rect 777 178 790 182
rect 796 179 820 183
rect 825 184 827 188
rect 707 170 721 174
rect 725 170 726 174
rect 777 173 780 178
rect 796 177 800 179
rect 766 169 780 173
rect 783 170 784 174
rect 788 170 789 174
rect 825 175 829 184
rect 854 182 858 194
rect 879 192 883 199
rect 887 197 888 201
rect 892 200 893 201
rect 892 197 904 200
rect 887 196 904 197
rect 900 193 904 196
rect 909 198 913 204
rect 923 201 927 208
rect 923 200 928 201
rect 909 195 916 198
rect 923 196 924 200
rect 931 200 935 221
rect 938 215 951 216
rect 938 211 941 215
rect 945 211 947 215
rect 938 210 951 211
rect 938 203 944 210
rect 954 204 958 221
rect 931 196 934 200
rect 938 196 939 200
rect 943 196 944 200
rect 948 196 949 200
rect 954 199 958 200
rect 923 195 928 196
rect 900 192 905 193
rect 868 186 874 191
rect 879 188 891 192
rect 895 188 896 192
rect 900 188 901 192
rect 868 184 870 186
rect 861 182 870 184
rect 900 187 905 188
rect 900 183 904 187
rect 861 178 874 182
rect 880 179 904 183
rect 854 177 858 178
rect 880 177 884 179
rect 796 172 800 173
rect 805 171 806 175
rect 810 171 829 175
rect 766 165 770 169
rect 783 165 789 170
rect 867 170 868 174
rect 872 170 873 174
rect 909 175 913 195
rect 923 187 927 195
rect 943 191 949 196
rect 930 187 931 191
rect 935 187 949 191
rect 955 190 959 192
rect 880 172 884 173
rect 889 171 890 175
rect 894 171 913 175
rect 917 184 927 187
rect 917 172 920 184
rect 867 165 873 170
rect 923 178 927 184
rect 923 177 928 178
rect 923 173 924 177
rect 928 173 935 176
rect 923 170 935 173
rect 939 174 943 187
rect 955 183 959 186
rect 946 179 950 183
rect 954 179 959 183
rect 946 178 959 179
rect 939 170 953 174
rect 957 170 958 174
rect 690 162 693 165
rect 689 161 693 162
rect 697 161 703 165
rect 707 161 771 165
rect 775 161 824 165
rect 828 161 855 165
rect 859 161 908 165
rect 912 161 925 165
rect 929 161 935 165
rect 939 161 963 165
rect 689 159 963 161
rect 670 158 963 159
rect 673 157 963 158
rect 673 156 692 157
rect 780 155 824 157
rect 780 151 786 155
rect 790 151 814 155
rect 818 151 824 155
rect 727 149 731 150
rect 671 131 700 136
rect 656 90 661 110
rect 727 108 731 145
rect 784 143 790 151
rect 784 139 785 143
rect 789 139 790 143
rect 795 143 799 144
rect 804 143 810 151
rect 804 139 805 143
rect 809 139 810 143
rect 815 143 820 146
rect 819 139 820 143
rect 795 136 799 139
rect 815 138 820 139
rect 795 132 812 136
rect 784 120 788 130
rect 792 125 797 129
rect 808 128 812 132
rect 792 117 798 121
rect 802 117 805 121
rect 792 111 796 117
rect 808 113 812 124
rect 779 108 796 111
rect 800 109 812 113
rect 816 133 832 138
rect 800 105 804 109
rect 816 108 820 133
rect 815 107 820 108
rect 784 101 785 105
rect 789 101 804 105
rect 807 103 815 105
rect 819 103 820 107
rect 807 101 820 103
rect 802 95 803 98
rect 780 94 803 95
rect 807 95 808 98
rect 807 94 814 95
rect 780 91 814 94
rect 818 91 824 95
rect 780 90 824 91
rect 656 87 824 90
rect 656 86 780 87
rect 978 82 981 237
rect 987 238 1348 241
rect 987 99 990 238
rect 1171 235 1176 238
rect 1277 235 1281 238
rect 1103 232 1352 235
rect 1103 227 1106 232
rect 1149 226 1152 232
rect 1203 226 1206 232
rect 1259 226 1262 232
rect 1313 226 1316 232
rect 1137 215 1140 223
rect 1137 211 1138 215
rect 1120 202 1123 205
rect 1137 189 1140 211
rect 1183 209 1186 222
rect 1183 206 1193 209
rect 1225 206 1228 210
rect 1237 212 1240 222
rect 1237 209 1256 212
rect 1285 212 1288 213
rect 1152 202 1154 205
rect 1174 202 1175 205
rect 1183 197 1186 206
rect 1150 194 1186 197
rect 1150 189 1153 194
rect 1183 189 1186 194
rect 1190 197 1193 206
rect 1204 202 1208 204
rect 1225 203 1229 206
rect 1204 201 1211 202
rect 1237 197 1240 209
rect 1287 208 1288 212
rect 1285 206 1288 208
rect 1261 202 1264 205
rect 1293 202 1296 222
rect 1319 215 1320 219
rect 1317 206 1320 215
rect 1347 211 1350 222
rect 1317 203 1318 206
rect 1336 202 1339 204
rect 1336 201 1342 202
rect 1293 197 1296 198
rect 1347 197 1350 207
rect 1204 194 1240 197
rect 1204 189 1207 194
rect 1237 189 1240 194
rect 1260 194 1296 197
rect 1260 189 1263 194
rect 1293 189 1296 194
rect 1314 194 1350 197
rect 1314 189 1317 194
rect 1347 189 1350 194
rect 1103 168 1106 185
rect 1166 168 1169 185
rect 1176 168 1179 171
rect 1220 168 1223 185
rect 1230 168 1233 171
rect 1276 168 1279 185
rect 1286 168 1289 171
rect 1330 168 1333 185
rect 1361 175 1366 307
rect 1372 306 1419 307
rect 1372 302 1378 306
rect 1382 302 1388 306
rect 1392 302 1419 306
rect 1391 296 1404 297
rect 1391 292 1399 296
rect 1403 292 1404 296
rect 1399 289 1404 292
rect 1376 284 1377 288
rect 1381 284 1396 288
rect 1403 285 1404 289
rect 1399 284 1404 285
rect 1374 277 1380 281
rect 1376 273 1380 277
rect 1376 272 1388 273
rect 1376 268 1380 272
rect 1384 268 1388 272
rect 1376 267 1388 268
rect 1392 272 1396 284
rect 1392 263 1396 268
rect 1400 271 1404 284
rect 1498 296 1504 312
rect 1520 311 1523 316
rect 1561 312 1575 318
rect 1567 308 1571 312
rect 1498 290 1514 296
rect 1567 295 1575 308
rect 1581 330 1585 331
rect 1581 311 1585 326
rect 1589 320 1593 336
rect 1598 337 1621 341
rect 1598 329 1602 337
rect 1617 334 1621 337
rect 1598 324 1602 325
rect 1606 332 1611 333
rect 1606 328 1607 332
rect 1617 330 1626 334
rect 1606 327 1611 328
rect 1606 320 1610 327
rect 1589 319 1610 320
rect 1589 316 1598 319
rect 1597 315 1598 316
rect 1602 316 1610 319
rect 1614 322 1618 323
rect 1602 315 1603 316
rect 1614 311 1618 318
rect 1581 309 1618 311
rect 1581 307 1594 309
rect 1598 307 1618 309
rect 1622 312 1626 330
rect 1622 307 1626 308
rect 1631 332 1655 344
rect 1635 328 1655 332
rect 1631 323 1655 328
rect 1631 319 1651 323
rect 1631 307 1655 319
rect 1660 343 1664 344
rect 1660 321 1664 339
rect 1668 342 1688 344
rect 1692 342 1705 344
rect 1668 340 1705 342
rect 1668 333 1672 340
rect 1683 335 1684 336
rect 1668 328 1672 329
rect 1676 332 1684 335
rect 1688 335 1689 336
rect 1688 332 1697 335
rect 1676 331 1697 332
rect 1676 324 1680 331
rect 1675 323 1680 324
rect 1660 317 1669 321
rect 1679 319 1680 323
rect 1675 318 1680 319
rect 1684 326 1688 327
rect 1665 314 1669 317
rect 1684 314 1688 322
rect 1665 310 1688 314
rect 1693 315 1697 331
rect 1701 325 1705 340
rect 1701 320 1705 321
rect 1711 343 1719 370
rect 1729 354 1745 357
rect 1715 339 1719 343
rect 1711 333 1725 339
rect 1742 335 1745 354
rect 1711 329 1721 333
rect 1730 334 1775 335
rect 1730 330 1733 334
rect 1737 331 1769 334
rect 1737 330 1738 331
rect 1768 330 1769 331
rect 1773 330 1775 334
rect 1711 325 1725 329
rect 1711 324 1737 325
rect 1711 320 1733 324
rect 1711 319 1737 320
rect 1740 323 1748 327
rect 1752 323 1767 327
rect 1693 311 1699 315
rect 1703 311 1704 315
rect 1533 291 1575 295
rect 1400 268 1449 271
rect 1400 264 1404 268
rect 1376 259 1377 263
rect 1381 259 1396 263
rect 1399 263 1404 264
rect 1403 259 1404 263
rect 1399 256 1404 259
rect 1387 251 1388 255
rect 1392 251 1393 255
rect 1403 252 1404 256
rect 1399 251 1404 252
rect 1387 246 1393 251
rect 1372 243 1378 246
rect 1373 242 1378 243
rect 1382 242 1414 246
rect 1373 240 1414 242
rect 1373 239 1426 240
rect 1372 238 1426 239
rect 1373 237 1426 238
rect 1373 233 1379 237
rect 1383 236 1426 237
rect 1383 233 1414 236
rect 1388 228 1394 233
rect 1388 224 1389 228
rect 1393 224 1394 228
rect 1400 227 1405 228
rect 1404 223 1405 227
rect 1400 220 1405 223
rect 1377 216 1378 220
rect 1382 216 1397 220
rect 1377 211 1389 212
rect 1377 207 1381 211
rect 1385 207 1389 211
rect 1377 206 1389 207
rect 1393 211 1397 216
rect 1404 216 1405 220
rect 1400 215 1405 216
rect 1377 202 1381 206
rect 1376 198 1381 202
rect 1393 195 1397 207
rect 1401 203 1405 215
rect 1401 199 1404 203
rect 1401 195 1405 199
rect 1377 191 1378 195
rect 1382 191 1397 195
rect 1400 194 1405 195
rect 1404 190 1405 194
rect 1400 187 1405 190
rect 1392 183 1400 187
rect 1404 183 1405 187
rect 1392 182 1405 183
rect 1373 175 1379 177
rect 1361 173 1379 175
rect 1383 173 1389 177
rect 1393 173 1408 177
rect 1361 172 1408 173
rect 1340 168 1343 171
rect 1361 168 1366 172
rect 999 165 1366 168
rect 1015 146 1018 165
rect 1098 163 1366 165
rect 1372 166 1408 172
rect 1049 158 1050 161
rect 1049 131 1052 158
rect 1060 148 1064 150
rect 1098 146 1101 163
rect 1109 154 1141 157
rect 1043 127 1046 130
rect 1050 128 1052 131
rect 1060 131 1064 142
rect 1060 121 1063 131
rect 1115 126 1118 129
rect 1060 117 1061 121
rect 1132 120 1135 142
rect 1138 130 1141 154
rect 1161 146 1164 163
rect 1171 160 1174 163
rect 1215 146 1218 163
rect 1225 160 1228 163
rect 1271 146 1274 163
rect 1281 160 1284 163
rect 1325 146 1328 163
rect 1335 160 1338 163
rect 1145 137 1148 142
rect 1178 137 1181 142
rect 1145 134 1181 137
rect 1138 127 1143 130
rect 1147 126 1149 129
rect 1169 126 1170 129
rect 1178 125 1181 134
rect 1199 137 1202 142
rect 1232 137 1235 142
rect 1199 134 1235 137
rect 1255 137 1258 142
rect 1288 137 1291 142
rect 1255 134 1291 137
rect 1309 137 1312 142
rect 1342 137 1345 142
rect 1309 134 1345 137
rect 1185 125 1188 134
rect 1199 129 1206 130
rect 1199 127 1203 129
rect 1220 125 1224 128
rect 1178 122 1188 125
rect 1060 109 1063 117
rect 1132 116 1133 120
rect 1132 108 1135 116
rect 1178 109 1181 122
rect 1220 121 1223 125
rect 1232 122 1235 134
rect 1288 133 1291 134
rect 1256 126 1259 129
rect 1232 119 1251 122
rect 1232 109 1235 119
rect 1280 123 1283 125
rect 1268 115 1271 121
rect 1282 119 1283 123
rect 1280 118 1283 119
rect 1245 112 1271 115
rect 1288 109 1291 129
rect 1312 125 1313 128
rect 1331 129 1337 130
rect 1331 127 1334 129
rect 1312 116 1315 125
rect 1342 124 1345 134
rect 1314 112 1315 116
rect 1342 109 1345 120
rect 1026 99 1029 105
rect 1098 99 1101 104
rect 1144 99 1147 105
rect 1198 99 1201 105
rect 1254 99 1257 105
rect 1308 99 1311 105
rect 986 96 1347 99
rect 1170 93 1175 96
rect 1276 93 1280 96
rect 1102 90 1351 93
rect 1102 85 1105 90
rect 1040 82 1044 83
rect 978 79 1045 82
rect 1148 84 1151 90
rect 1202 84 1205 90
rect 1258 84 1261 90
rect 1312 84 1315 90
rect 622 53 626 78
rect 904 73 908 74
rect 682 69 908 73
rect 904 65 908 69
rect 904 63 1015 65
rect 1020 63 1023 65
rect 904 60 1023 63
rect 622 52 745 53
rect 622 51 991 52
rect 622 48 1007 51
rect 1020 44 1023 60
rect 1015 41 1023 44
rect 524 34 527 38
rect 531 34 538 38
rect 585 34 990 38
rect 517 30 521 34
rect 517 26 529 30
rect 509 24 514 25
rect 438 18 453 22
rect 457 18 458 22
rect 509 20 510 24
rect 514 20 521 23
rect 509 17 521 20
rect 525 22 529 26
rect 533 28 538 34
rect 533 25 546 28
rect 551 26 999 29
rect 1040 27 1044 79
rect 1136 73 1139 81
rect 1136 69 1137 73
rect 1119 60 1122 63
rect 1093 48 1096 49
rect 1063 45 1096 48
rect 1136 47 1139 69
rect 1182 67 1185 80
rect 1182 64 1192 67
rect 1224 64 1227 68
rect 1236 70 1239 80
rect 1236 67 1255 70
rect 1284 70 1287 71
rect 1151 60 1153 63
rect 1173 60 1174 63
rect 1182 55 1185 64
rect 1149 52 1185 55
rect 1149 47 1152 52
rect 1182 47 1185 52
rect 1189 55 1192 64
rect 1203 60 1207 62
rect 1224 61 1228 64
rect 1203 59 1210 60
rect 1236 55 1239 67
rect 1286 66 1287 70
rect 1284 64 1287 66
rect 1260 60 1263 63
rect 1292 60 1295 80
rect 1318 73 1319 77
rect 1316 64 1319 73
rect 1346 69 1349 80
rect 1316 61 1317 64
rect 1335 60 1338 62
rect 1335 59 1341 60
rect 1292 55 1295 56
rect 1346 55 1349 65
rect 1203 52 1239 55
rect 1203 47 1206 52
rect 1236 47 1239 52
rect 1259 52 1295 55
rect 1259 47 1262 52
rect 1292 47 1295 52
rect 1313 52 1349 55
rect 1313 47 1316 52
rect 1346 47 1349 52
rect 1093 41 1096 45
rect 1058 37 1096 41
rect 1058 34 1061 37
rect 1088 29 1091 32
rect 1096 29 1097 32
rect 1088 27 1097 29
rect 1040 23 1097 27
rect 1102 24 1105 43
rect 1165 24 1168 43
rect 1175 24 1178 29
rect 1219 24 1222 43
rect 1229 24 1232 29
rect 1275 24 1278 43
rect 1285 24 1288 29
rect 1329 24 1332 43
rect 1339 24 1342 29
rect 1360 24 1365 163
rect 1372 162 1378 166
rect 1382 162 1388 166
rect 1392 162 1408 166
rect 1391 156 1404 157
rect 1391 152 1399 156
rect 1403 152 1404 156
rect 1399 149 1404 152
rect 1376 144 1377 148
rect 1381 144 1396 148
rect 1403 145 1404 149
rect 1399 144 1404 145
rect 1376 133 1380 141
rect 1376 132 1388 133
rect 1376 128 1380 132
rect 1384 128 1388 132
rect 1376 127 1388 128
rect 1392 132 1396 144
rect 1392 123 1396 128
rect 1400 136 1404 144
rect 1400 132 1403 136
rect 1400 124 1404 132
rect 1376 119 1377 123
rect 1381 119 1396 123
rect 1399 123 1404 124
rect 1403 119 1404 123
rect 1399 116 1404 119
rect 1387 111 1388 115
rect 1392 111 1393 115
rect 1403 112 1404 116
rect 1399 111 1404 112
rect 1387 106 1393 111
rect 1411 106 1414 233
rect 1372 102 1378 106
rect 1382 102 1414 106
rect 1372 98 1414 102
rect 1395 70 1399 91
rect 1437 72 1441 268
rect 525 18 540 22
rect 544 18 545 22
rect 1100 21 1365 24
rect 1379 67 1399 70
rect 1379 23 1383 67
rect 1438 62 1441 72
rect 1498 137 1504 290
rect 1533 261 1538 291
rect 1514 257 1538 261
rect 1514 208 1518 257
rect 1533 256 1538 257
rect 1567 281 1575 291
rect 1631 303 1654 307
rect 1658 303 1661 307
rect 1665 303 1666 307
rect 1612 282 1626 283
rect 1567 277 1571 281
rect 1587 278 1588 282
rect 1592 278 1608 282
rect 1612 278 1613 282
rect 1617 278 1626 282
rect 1567 269 1575 277
rect 1567 268 1584 269
rect 1567 264 1580 268
rect 1567 263 1584 264
rect 1588 268 1594 275
rect 1604 274 1608 278
rect 1620 274 1621 278
rect 1625 274 1626 278
rect 1604 270 1607 274
rect 1611 270 1613 274
rect 1620 271 1626 274
rect 1588 266 1601 268
rect 1515 203 1518 208
rect 1541 193 1545 229
rect 1516 189 1545 193
rect 1553 149 1556 239
rect 1560 208 1563 226
rect 1567 228 1575 263
rect 1588 262 1592 266
rect 1596 262 1601 266
rect 1609 257 1613 270
rect 1631 264 1655 303
rect 1673 297 1677 310
rect 1711 305 1725 319
rect 1740 314 1744 323
rect 1755 317 1759 320
rect 1732 310 1733 314
rect 1737 310 1744 314
rect 1763 319 1767 323
rect 1771 322 1775 330
rect 1781 333 1789 339
rect 1785 329 1789 333
rect 1781 323 1789 329
rect 1778 322 1789 323
rect 1763 315 1775 319
rect 1782 318 1789 322
rect 1778 317 1789 318
rect 1747 307 1751 312
rect 1755 311 1759 313
rect 1755 307 1768 311
rect 1685 301 1690 305
rect 1694 301 1698 305
rect 1711 304 1721 305
rect 1685 299 1698 301
rect 1660 289 1666 296
rect 1673 293 1675 297
rect 1679 293 1682 297
rect 1678 289 1682 293
rect 1692 292 1698 299
rect 1702 303 1721 304
rect 1706 301 1721 303
rect 1725 304 1737 305
rect 1725 301 1733 304
rect 1706 300 1733 301
rect 1706 299 1737 300
rect 1746 299 1756 303
rect 1702 298 1725 299
rect 1711 295 1725 298
rect 1711 290 1719 295
rect 1765 294 1768 307
rect 1771 304 1775 315
rect 1771 299 1775 300
rect 1781 295 1789 317
rect 1660 285 1669 289
rect 1673 285 1674 289
rect 1678 285 1694 289
rect 1698 285 1699 289
rect 1715 286 1719 290
rect 1660 284 1674 285
rect 1670 279 1673 284
rect 1670 276 1687 279
rect 1620 260 1621 264
rect 1625 260 1628 264
rect 1632 260 1655 264
rect 1582 252 1583 256
rect 1587 252 1593 256
rect 1567 224 1571 228
rect 1567 211 1575 224
rect 1581 246 1585 247
rect 1581 227 1585 242
rect 1589 236 1593 252
rect 1598 253 1621 257
rect 1598 245 1602 253
rect 1617 250 1621 253
rect 1598 240 1602 241
rect 1606 248 1611 249
rect 1606 244 1607 248
rect 1617 246 1626 250
rect 1606 243 1611 244
rect 1606 236 1610 243
rect 1589 235 1610 236
rect 1589 232 1598 235
rect 1597 231 1598 232
rect 1602 232 1610 235
rect 1614 238 1618 239
rect 1602 231 1603 232
rect 1614 227 1618 234
rect 1581 223 1618 227
rect 1622 228 1626 246
rect 1622 223 1626 224
rect 1631 248 1655 260
rect 1635 244 1655 248
rect 1631 241 1655 244
rect 1711 269 1719 286
rect 1631 240 1672 241
rect 1631 236 1651 240
rect 1655 237 1672 240
rect 1676 237 1677 241
rect 1684 238 1687 242
rect 1691 238 1698 242
rect 1693 237 1698 238
rect 1631 226 1655 236
rect 1605 220 1608 223
rect 1582 216 1597 219
rect 1631 222 1651 226
rect 1631 218 1655 222
rect 1660 230 1661 234
rect 1665 230 1666 234
rect 1697 233 1698 237
rect 1660 228 1666 230
rect 1660 224 1661 228
rect 1665 227 1666 228
rect 1676 231 1689 232
rect 1680 227 1689 231
rect 1693 229 1698 233
rect 1702 240 1706 241
rect 1665 224 1673 227
rect 1676 226 1689 227
rect 1702 226 1706 236
rect 1660 221 1673 224
rect 1685 222 1706 226
rect 1711 222 1725 269
rect 1748 256 1775 257
rect 1748 254 1772 256
rect 1676 221 1680 222
rect 1631 217 1676 218
rect 1594 213 1597 216
rect 1631 214 1680 217
rect 1685 218 1689 222
rect 1715 218 1725 222
rect 1567 207 1571 211
rect 1567 201 1575 207
rect 1580 212 1618 213
rect 1580 208 1583 212
rect 1587 209 1606 212
rect 1587 208 1588 209
rect 1605 208 1606 209
rect 1610 209 1618 212
rect 1631 212 1655 214
rect 1685 213 1689 214
rect 1631 211 1651 212
rect 1610 208 1611 209
rect 1580 201 1586 208
rect 1635 208 1651 211
rect 1700 211 1706 218
rect 1675 210 1676 211
rect 1635 207 1655 208
rect 1597 205 1601 206
rect 1631 205 1655 207
rect 1668 207 1676 210
rect 1680 210 1681 211
rect 1698 210 1699 211
rect 1680 207 1689 210
rect 1668 206 1689 207
rect 1693 207 1699 210
rect 1703 207 1706 211
rect 1693 206 1706 207
rect 1711 212 1725 218
rect 1715 208 1725 212
rect 1711 205 1725 208
rect 1567 197 1571 201
rect 1597 197 1601 201
rect 1606 202 1655 205
rect 1610 201 1655 202
rect 1606 197 1610 198
rect 1567 173 1575 197
rect 1580 193 1601 197
rect 1613 195 1626 198
rect 1580 183 1584 193
rect 1597 192 1610 193
rect 1613 192 1621 195
rect 1580 178 1584 179
rect 1588 186 1593 190
rect 1597 188 1606 192
rect 1597 187 1610 188
rect 1620 191 1621 192
rect 1625 191 1626 195
rect 1620 189 1626 191
rect 1588 182 1589 186
rect 1620 185 1621 189
rect 1625 185 1626 189
rect 1631 197 1655 201
rect 1635 193 1655 197
rect 1631 183 1655 193
rect 1715 191 1725 205
rect 1715 188 1717 191
rect 1588 181 1593 182
rect 1588 177 1596 181
rect 1600 177 1602 181
rect 1609 178 1610 182
rect 1614 179 1631 182
rect 1635 179 1655 183
rect 1614 178 1655 179
rect 1631 176 1655 178
rect 1786 176 1790 295
rect 1631 175 1790 176
rect 1631 173 1791 175
rect 1511 148 1556 149
rect 1515 145 1556 148
rect 1569 145 1574 173
rect 1647 172 1791 173
rect 1766 171 1791 172
rect 1569 144 1695 145
rect 1569 139 1690 144
rect 1715 143 1720 148
rect 1697 138 1720 143
rect 1692 137 1720 138
rect 1498 119 1502 137
rect 1715 136 1720 137
rect 1715 133 1719 136
rect 1526 128 1547 132
rect 1509 119 1522 120
rect 1498 118 1651 119
rect 1715 118 1720 133
rect 1726 121 1729 157
rect 1498 115 1657 118
rect 1392 59 1442 62
rect 182 7 188 13
rect 187 0 188 7
rect 325 8 331 12
rect 335 8 341 12
rect 345 8 369 12
rect 418 8 424 12
rect 428 8 434 12
rect 438 8 462 12
rect 319 7 462 8
rect 505 8 511 12
rect 515 8 521 12
rect 525 8 549 12
rect 505 7 549 8
rect 319 5 549 7
rect 325 4 369 5
rect 418 4 549 5
rect 981 5 1048 8
rect 1392 7 1396 59
rect 1419 19 1441 23
rect -14 -8 -6 -4
rect 981 -8 985 5
rect -14 -13 985 -8
rect 1007 0 1010 1
rect 1393 0 1396 7
rect 1007 -4 1398 0
rect -14 -82 -6 -13
rect 983 -26 998 -22
rect 44 -48 485 -44
rect 44 -70 48 -48
rect 126 -57 127 -54
rect 342 -57 535 -56
rect 541 -57 585 -55
rect 126 -58 585 -57
rect 634 -58 678 -55
rect 721 -56 765 -55
rect 721 -58 773 -56
rect 121 -59 773 -58
rect 121 -61 547 -59
rect 121 -65 145 -61
rect 149 -65 155 -61
rect 159 -65 232 -61
rect 236 -65 242 -61
rect 246 -65 325 -61
rect 329 -65 335 -61
rect 339 -62 547 -61
rect 339 -65 345 -62
rect 541 -63 547 -62
rect 551 -63 557 -59
rect 561 -62 640 -59
rect 561 -63 585 -62
rect 634 -63 640 -62
rect 644 -63 650 -59
rect 654 -62 727 -59
rect 654 -63 678 -62
rect 721 -63 727 -62
rect 731 -63 737 -59
rect 741 -62 773 -59
rect 741 -63 765 -62
rect 125 -75 126 -71
rect 130 -75 145 -71
rect 82 -82 121 -79
rect 125 -82 137 -78
rect -14 -84 46 -82
rect 82 -84 85 -82
rect -14 -87 85 -84
rect 132 -87 137 -82
rect 141 -79 145 -75
rect 149 -73 161 -70
rect 149 -76 156 -73
rect 160 -77 161 -73
rect 212 -75 213 -71
rect 217 -75 232 -71
rect 156 -78 161 -77
rect 141 -83 153 -79
rect 149 -87 153 -83
rect -14 -89 46 -87
rect 132 -91 139 -87
rect 143 -91 146 -87
rect 125 -104 129 -95
rect 133 -99 138 -95
rect 149 -102 153 -91
rect 157 -92 161 -78
rect 213 -82 224 -78
rect 219 -87 224 -82
rect 228 -79 232 -75
rect 236 -73 248 -70
rect 236 -76 243 -73
rect 247 -77 248 -73
rect 305 -75 306 -71
rect 310 -75 325 -71
rect 243 -78 248 -77
rect 228 -83 240 -79
rect 236 -87 240 -83
rect 219 -91 226 -87
rect 230 -91 233 -87
rect 157 -95 186 -92
rect 157 -96 161 -95
rect 118 -108 129 -104
rect 136 -104 153 -102
rect 140 -106 153 -104
rect 156 -97 161 -96
rect 160 -101 161 -97
rect 156 -104 161 -101
rect 136 -111 140 -108
rect 160 -108 161 -104
rect 156 -109 161 -108
rect 125 -115 126 -111
rect 130 -115 131 -111
rect 125 -121 131 -115
rect 136 -116 140 -115
rect 145 -113 146 -109
rect 150 -113 151 -109
rect 145 -121 151 -113
rect 121 -125 155 -121
rect 159 -125 165 -121
rect 121 -129 165 -125
rect -37 -136 24 -134
rect 122 -136 126 -129
rect 182 -131 186 -95
rect 212 -105 216 -95
rect 220 -99 225 -95
rect 236 -102 240 -91
rect 244 -96 248 -78
rect 306 -82 317 -78
rect 312 -87 317 -82
rect 321 -79 325 -75
rect 329 -73 341 -70
rect 545 -71 557 -68
rect 329 -76 336 -73
rect 340 -77 341 -73
rect 354 -77 423 -73
rect 429 -77 526 -73
rect 531 -77 532 -73
rect 545 -75 546 -71
rect 550 -74 557 -71
rect 561 -73 576 -69
rect 580 -73 581 -69
rect 638 -71 650 -68
rect 545 -76 550 -75
rect 336 -78 341 -77
rect 321 -83 333 -79
rect 329 -87 333 -83
rect 312 -91 319 -87
rect 323 -91 326 -87
rect 209 -108 216 -105
rect 223 -104 240 -102
rect 227 -106 240 -104
rect 243 -97 248 -96
rect 247 -101 248 -97
rect 243 -104 248 -101
rect 223 -111 227 -108
rect 247 -106 248 -104
rect 247 -108 254 -106
rect 243 -109 254 -108
rect 305 -105 309 -95
rect 313 -99 318 -95
rect 329 -102 333 -91
rect 337 -83 341 -78
rect 337 -86 431 -83
rect 337 -96 341 -86
rect 545 -83 549 -76
rect 561 -77 565 -73
rect 638 -75 639 -71
rect 643 -74 650 -71
rect 654 -73 669 -69
rect 673 -73 674 -69
rect 725 -71 737 -68
rect 638 -76 643 -75
rect 489 -87 549 -83
rect 302 -108 309 -105
rect 316 -104 333 -102
rect 320 -106 333 -104
rect 336 -97 341 -96
rect 340 -101 341 -97
rect 354 -99 411 -96
rect 545 -94 549 -87
rect 553 -81 565 -77
rect 569 -79 580 -76
rect 553 -85 557 -81
rect 569 -85 574 -79
rect 560 -89 563 -85
rect 567 -89 574 -85
rect 638 -87 642 -76
rect 654 -77 658 -73
rect 725 -75 726 -71
rect 730 -74 737 -71
rect 741 -73 756 -69
rect 760 -73 761 -69
rect 725 -76 730 -75
rect 545 -95 550 -94
rect 417 -99 527 -96
rect 545 -99 546 -95
rect 336 -104 341 -101
rect 545 -102 550 -99
rect 212 -115 213 -111
rect 217 -115 218 -111
rect 212 -121 218 -115
rect 223 -116 227 -115
rect 232 -113 233 -109
rect 237 -113 238 -109
rect 316 -111 320 -108
rect 340 -108 341 -104
rect 336 -109 341 -108
rect 232 -121 238 -113
rect 305 -115 306 -111
rect 310 -115 311 -111
rect 305 -121 311 -115
rect 316 -116 320 -115
rect 325 -113 326 -109
rect 330 -113 331 -109
rect 491 -109 513 -105
rect 545 -106 546 -102
rect 553 -100 557 -89
rect 615 -90 642 -87
rect 568 -97 573 -93
rect 553 -102 570 -100
rect 553 -104 566 -102
rect 545 -107 550 -106
rect 577 -103 581 -93
rect 615 -102 619 -90
rect 577 -106 584 -103
rect 325 -121 331 -113
rect 392 -114 396 -110
rect 555 -111 556 -107
rect 560 -111 561 -107
rect 354 -117 528 -114
rect 555 -119 561 -111
rect 566 -109 570 -106
rect 638 -94 642 -90
rect 646 -81 658 -77
rect 662 -77 676 -76
rect 662 -79 673 -77
rect 646 -85 650 -81
rect 662 -85 667 -79
rect 653 -89 656 -85
rect 660 -89 667 -85
rect 638 -95 643 -94
rect 638 -99 639 -95
rect 638 -102 643 -99
rect 638 -106 639 -102
rect 646 -100 650 -89
rect 725 -90 729 -76
rect 741 -77 745 -73
rect 661 -97 666 -93
rect 646 -102 663 -100
rect 646 -104 659 -102
rect 638 -107 643 -106
rect 670 -103 674 -93
rect 703 -94 729 -90
rect 733 -81 745 -77
rect 749 -77 763 -76
rect 749 -79 760 -77
rect 733 -85 737 -81
rect 749 -85 754 -79
rect 1007 -78 1010 -4
rect 1023 -11 1056 -7
rect 1052 -14 1056 -11
rect 1109 -11 1112 -4
rect 1052 -18 1053 -14
rect 1021 -26 1131 -22
rect 1018 -27 1131 -26
rect 1407 -35 1412 -33
rect 1104 -38 1412 -35
rect 1021 -59 1387 -56
rect 1037 -78 1040 -59
rect 1082 -76 1086 -74
rect 764 -81 1011 -78
rect 740 -89 743 -85
rect 747 -89 754 -85
rect 670 -106 677 -103
rect 689 -104 690 -100
rect 566 -114 570 -113
rect 575 -113 576 -109
rect 580 -113 581 -109
rect 575 -119 581 -113
rect 648 -111 649 -107
rect 653 -111 654 -107
rect 648 -119 654 -111
rect 659 -109 663 -106
rect 659 -114 663 -113
rect 668 -113 669 -109
rect 673 -113 674 -109
rect 668 -119 674 -113
rect 208 -125 242 -121
rect 246 -125 252 -121
rect 208 -126 252 -125
rect 301 -125 335 -121
rect 339 -125 345 -121
rect 208 -129 235 -126
rect 301 -129 345 -125
rect 541 -123 547 -119
rect 551 -123 585 -119
rect 634 -123 640 -119
rect 644 -123 678 -119
rect 541 -127 585 -123
rect 210 -136 214 -129
rect 247 -133 280 -130
rect 301 -136 305 -129
rect 577 -131 581 -127
rect 596 -128 626 -125
rect 634 -127 678 -123
rect 689 -124 693 -104
rect 535 -132 639 -131
rect 535 -134 661 -132
rect 670 -134 674 -127
rect 703 -125 707 -94
rect 725 -95 730 -94
rect 725 -99 726 -95
rect 713 -124 717 -104
rect 725 -102 730 -99
rect 725 -106 726 -102
rect 733 -100 737 -89
rect 748 -97 753 -93
rect 733 -102 750 -100
rect 733 -104 746 -102
rect 725 -107 730 -106
rect 757 -102 761 -93
rect 994 -95 1039 -92
rect 1082 -93 1086 -82
rect 1065 -97 1068 -94
rect 757 -106 765 -102
rect 1082 -103 1085 -93
rect 1109 -96 1112 -72
rect 1120 -78 1123 -59
rect 1183 -78 1186 -59
rect 1193 -64 1196 -59
rect 1237 -78 1240 -59
rect 1247 -64 1250 -59
rect 1293 -78 1296 -59
rect 1303 -64 1306 -59
rect 1347 -78 1350 -59
rect 1357 -64 1360 -59
rect 1109 -99 1133 -96
rect 1137 -98 1140 -95
rect 735 -111 736 -107
rect 740 -111 741 -107
rect 735 -119 741 -111
rect 746 -109 750 -106
rect 1082 -107 1083 -103
rect 1154 -104 1157 -82
rect 1167 -87 1170 -82
rect 1200 -87 1203 -82
rect 1167 -90 1203 -87
rect 1169 -98 1171 -95
rect 1191 -98 1192 -95
rect 1200 -99 1203 -90
rect 1221 -87 1224 -82
rect 1254 -87 1257 -82
rect 1221 -90 1257 -87
rect 1277 -87 1280 -82
rect 1310 -87 1313 -82
rect 1277 -90 1313 -87
rect 1331 -87 1334 -82
rect 1364 -87 1367 -82
rect 1331 -90 1367 -87
rect 1207 -99 1210 -90
rect 1221 -95 1228 -94
rect 1221 -97 1225 -95
rect 1242 -99 1246 -96
rect 1200 -102 1210 -99
rect 746 -114 750 -113
rect 755 -113 756 -109
rect 760 -113 761 -109
rect 755 -119 761 -113
rect 1082 -115 1085 -107
rect 1154 -108 1155 -104
rect 1154 -116 1157 -108
rect 1200 -115 1203 -102
rect 1242 -103 1245 -99
rect 1254 -102 1257 -90
rect 1310 -91 1313 -90
rect 1278 -98 1281 -95
rect 1254 -105 1273 -102
rect 1254 -115 1257 -105
rect 1302 -101 1305 -99
rect 1290 -109 1293 -103
rect 1304 -105 1305 -101
rect 1302 -106 1305 -105
rect 1267 -112 1293 -109
rect 1310 -115 1313 -95
rect 1334 -99 1335 -96
rect 1353 -95 1359 -94
rect 1353 -97 1356 -95
rect 1334 -108 1337 -99
rect 1364 -100 1367 -90
rect 1336 -112 1337 -108
rect 1364 -115 1367 -104
rect 721 -123 727 -119
rect 731 -123 765 -119
rect 721 -127 765 -123
rect 1048 -125 1051 -119
rect 1120 -125 1123 -120
rect 1166 -125 1169 -119
rect 1220 -125 1223 -119
rect 1276 -125 1279 -119
rect 1330 -125 1333 -119
rect 759 -134 763 -127
rect 1012 -128 1369 -125
rect 1012 -129 1027 -128
rect 773 -134 975 -131
rect 317 -135 975 -134
rect 317 -136 705 -135
rect -37 -137 240 -136
rect 253 -137 705 -136
rect -37 -138 705 -137
rect -37 -140 378 -138
rect -37 -144 49 -140
rect 53 -144 63 -140
rect 67 -144 77 -140
rect 81 -143 160 -140
rect 81 -144 144 -143
rect -37 -146 24 -144
rect 33 -145 48 -144
rect 13 -255 17 -146
rect 47 -164 51 -157
rect 47 -165 52 -164
rect 47 -169 48 -165
rect 55 -165 59 -144
rect 62 -150 75 -149
rect 62 -154 65 -150
rect 69 -154 71 -150
rect 62 -155 75 -154
rect 62 -162 68 -155
rect 78 -161 82 -144
rect 148 -144 160 -143
rect 164 -143 244 -140
rect 164 -144 228 -143
rect 125 -155 137 -149
rect 144 -150 148 -147
rect 232 -144 244 -143
rect 248 -144 281 -140
rect 285 -144 295 -140
rect 299 -144 309 -140
rect 313 -142 378 -140
rect 382 -142 392 -138
rect 396 -142 406 -138
rect 410 -141 489 -138
rect 410 -142 473 -141
rect 313 -144 348 -142
rect 158 -153 180 -149
rect 184 -153 185 -149
rect 209 -150 221 -149
rect 158 -154 162 -153
rect 144 -155 148 -154
rect 125 -158 130 -155
rect 125 -159 126 -158
rect 55 -169 58 -165
rect 62 -169 63 -165
rect 67 -169 68 -165
rect 72 -169 73 -165
rect 78 -166 82 -165
rect 117 -162 126 -159
rect 151 -158 162 -154
rect 209 -154 214 -150
rect 218 -154 221 -150
rect 209 -155 221 -154
rect 228 -150 232 -147
rect 242 -153 264 -149
rect 268 -153 269 -149
rect 242 -154 246 -153
rect 228 -155 232 -154
rect 151 -162 155 -158
rect 169 -161 170 -157
rect 174 -161 185 -157
rect 47 -170 52 -169
rect 47 -178 51 -170
rect 67 -174 73 -169
rect 54 -178 55 -174
rect 59 -178 73 -174
rect 79 -176 83 -173
rect 117 -176 120 -162
rect 125 -163 130 -162
rect 134 -164 155 -162
rect 47 -187 51 -182
rect 47 -188 52 -187
rect 47 -192 48 -188
rect 52 -192 59 -189
rect 47 -195 59 -192
rect 63 -191 67 -178
rect 126 -168 134 -167
rect 138 -166 155 -164
rect 126 -171 138 -168
rect 79 -182 83 -180
rect 70 -186 74 -182
rect 78 -186 83 -182
rect 70 -187 83 -186
rect 126 -183 130 -171
rect 151 -173 155 -166
rect 159 -168 160 -164
rect 164 -165 165 -164
rect 164 -168 176 -165
rect 159 -169 176 -168
rect 172 -172 176 -169
rect 172 -173 177 -172
rect 140 -179 146 -174
rect 151 -177 163 -173
rect 167 -177 168 -173
rect 172 -177 173 -173
rect 140 -181 142 -179
rect 133 -183 142 -181
rect 172 -178 177 -177
rect 181 -177 185 -161
rect 209 -158 214 -155
rect 209 -162 210 -158
rect 235 -158 246 -154
rect 235 -162 239 -158
rect 253 -161 254 -157
rect 258 -161 269 -157
rect 209 -163 214 -162
rect 218 -164 239 -162
rect 210 -168 218 -167
rect 222 -166 239 -164
rect 210 -171 222 -168
rect 172 -182 176 -178
rect 133 -187 146 -183
rect 152 -186 176 -182
rect 181 -181 183 -177
rect 126 -188 130 -187
rect 152 -188 156 -186
rect 63 -195 77 -191
rect 81 -195 82 -191
rect 139 -195 140 -191
rect 144 -195 145 -191
rect 181 -190 185 -181
rect 210 -183 214 -171
rect 235 -173 239 -166
rect 243 -168 244 -164
rect 248 -165 249 -164
rect 248 -168 260 -165
rect 243 -169 260 -168
rect 256 -172 260 -169
rect 265 -170 269 -161
rect 279 -164 283 -157
rect 279 -165 284 -164
rect 279 -169 280 -165
rect 287 -165 291 -144
rect 294 -150 303 -149
rect 294 -154 297 -150
rect 301 -153 303 -150
rect 301 -154 307 -153
rect 294 -155 307 -154
rect 294 -162 300 -155
rect 310 -161 314 -144
rect 321 -161 339 -158
rect 287 -169 290 -165
rect 294 -169 295 -165
rect 299 -169 300 -165
rect 304 -169 305 -165
rect 310 -166 314 -165
rect 256 -173 261 -172
rect 224 -179 230 -174
rect 235 -177 247 -173
rect 251 -177 252 -173
rect 256 -177 257 -173
rect 224 -181 226 -179
rect 217 -183 226 -181
rect 256 -178 261 -177
rect 265 -173 272 -170
rect 279 -170 284 -169
rect 256 -182 260 -178
rect 217 -187 230 -183
rect 236 -186 260 -182
rect 210 -188 214 -187
rect 236 -188 240 -186
rect 152 -193 156 -192
rect 161 -194 162 -190
rect 166 -194 185 -190
rect 139 -200 145 -195
rect 223 -195 224 -191
rect 228 -195 229 -191
rect 265 -190 269 -173
rect 279 -178 283 -170
rect 299 -174 305 -169
rect 286 -178 287 -174
rect 291 -178 305 -174
rect 311 -175 315 -173
rect 236 -193 240 -192
rect 245 -194 246 -190
rect 250 -194 269 -190
rect 273 -181 283 -178
rect 273 -193 276 -181
rect 223 -200 229 -195
rect 279 -187 283 -181
rect 279 -188 284 -187
rect 279 -192 280 -188
rect 284 -192 291 -189
rect 279 -195 291 -192
rect 295 -191 299 -178
rect 311 -182 315 -179
rect 302 -186 306 -182
rect 310 -186 315 -182
rect 302 -187 315 -186
rect 295 -195 309 -191
rect 313 -195 314 -191
rect 46 -204 49 -200
rect 53 -204 59 -200
rect 63 -204 127 -200
rect 131 -204 180 -200
rect 184 -204 211 -200
rect 215 -204 264 -200
rect 268 -204 281 -200
rect 285 -204 291 -200
rect 295 -201 319 -200
rect 295 -204 313 -201
rect 32 -207 313 -204
rect 32 -208 319 -207
rect 136 -210 180 -208
rect 136 -214 142 -210
rect 146 -214 170 -210
rect 174 -214 180 -210
rect 140 -222 146 -214
rect 140 -226 141 -222
rect 145 -226 146 -222
rect 151 -222 155 -221
rect 160 -222 166 -214
rect 160 -226 161 -222
rect 165 -226 166 -222
rect 171 -222 176 -219
rect 334 -218 338 -161
rect 307 -221 339 -218
rect 175 -226 176 -222
rect 151 -229 155 -226
rect 171 -227 176 -226
rect 151 -233 168 -229
rect 140 -245 144 -235
rect 148 -240 153 -236
rect 164 -237 168 -233
rect 148 -248 154 -244
rect 158 -248 161 -244
rect 12 -275 17 -255
rect 148 -254 152 -248
rect 164 -252 168 -241
rect 135 -257 152 -254
rect 156 -256 168 -252
rect 172 -231 333 -227
rect 156 -260 160 -256
rect 172 -257 176 -231
rect 342 -253 346 -144
rect 376 -162 380 -155
rect 376 -163 381 -162
rect 376 -167 377 -163
rect 384 -163 388 -142
rect 391 -148 404 -147
rect 391 -152 394 -148
rect 398 -152 400 -148
rect 391 -153 404 -152
rect 391 -160 397 -153
rect 407 -159 411 -142
rect 477 -142 489 -141
rect 493 -141 573 -138
rect 493 -142 557 -141
rect 454 -153 466 -147
rect 473 -148 477 -145
rect 561 -142 573 -141
rect 577 -142 610 -138
rect 614 -142 624 -138
rect 628 -142 638 -138
rect 642 -139 705 -138
rect 709 -139 719 -135
rect 723 -139 733 -135
rect 737 -138 816 -135
rect 737 -139 800 -138
rect 642 -142 678 -139
rect 487 -151 509 -147
rect 513 -151 514 -147
rect 529 -148 550 -147
rect 487 -152 491 -151
rect 473 -153 477 -152
rect 454 -156 459 -153
rect 454 -157 455 -156
rect 384 -167 387 -163
rect 391 -167 392 -163
rect 396 -167 397 -163
rect 401 -167 402 -163
rect 407 -164 411 -163
rect 446 -160 455 -157
rect 480 -156 491 -152
rect 529 -152 543 -148
rect 547 -152 550 -148
rect 529 -153 550 -152
rect 557 -148 561 -145
rect 571 -151 593 -147
rect 597 -151 598 -147
rect 571 -152 575 -151
rect 557 -153 561 -152
rect 480 -160 484 -156
rect 498 -159 499 -155
rect 503 -159 514 -155
rect 376 -168 381 -167
rect 376 -176 380 -168
rect 396 -172 402 -167
rect 383 -176 384 -172
rect 388 -176 402 -172
rect 408 -174 412 -171
rect 446 -174 449 -160
rect 454 -161 459 -160
rect 463 -162 484 -160
rect 376 -185 380 -180
rect 376 -186 381 -185
rect 376 -190 377 -186
rect 381 -190 388 -187
rect 376 -193 388 -190
rect 392 -189 396 -176
rect 455 -166 463 -165
rect 467 -164 484 -162
rect 455 -169 467 -166
rect 408 -180 412 -178
rect 399 -184 403 -180
rect 407 -184 412 -180
rect 399 -185 412 -184
rect 455 -181 459 -169
rect 480 -171 484 -164
rect 488 -166 489 -162
rect 493 -163 494 -162
rect 493 -166 505 -163
rect 488 -167 505 -166
rect 501 -170 505 -167
rect 501 -171 506 -170
rect 469 -177 475 -172
rect 480 -175 492 -171
rect 496 -175 497 -171
rect 501 -175 502 -171
rect 469 -179 471 -177
rect 462 -181 471 -179
rect 501 -176 506 -175
rect 510 -175 514 -159
rect 538 -156 543 -153
rect 538 -160 539 -156
rect 564 -156 575 -152
rect 564 -160 568 -156
rect 582 -159 583 -155
rect 587 -159 600 -155
rect 538 -161 543 -160
rect 547 -162 568 -160
rect 539 -166 547 -165
rect 551 -164 568 -162
rect 539 -169 551 -166
rect 501 -180 505 -176
rect 462 -185 475 -181
rect 481 -184 505 -180
rect 510 -179 512 -175
rect 455 -186 459 -185
rect 481 -186 485 -184
rect 392 -193 406 -189
rect 410 -193 411 -189
rect 468 -193 469 -189
rect 473 -193 474 -189
rect 510 -188 514 -179
rect 539 -181 543 -169
rect 564 -171 568 -164
rect 572 -166 573 -162
rect 577 -163 578 -162
rect 577 -166 589 -163
rect 572 -167 589 -166
rect 585 -170 589 -167
rect 585 -171 590 -170
rect 553 -177 559 -172
rect 564 -175 576 -171
rect 580 -175 581 -171
rect 585 -175 586 -171
rect 553 -179 555 -177
rect 546 -181 555 -179
rect 585 -176 590 -175
rect 585 -180 589 -176
rect 546 -185 559 -181
rect 565 -184 589 -180
rect 539 -186 543 -185
rect 565 -186 569 -184
rect 481 -191 485 -190
rect 490 -192 491 -188
rect 495 -192 514 -188
rect 468 -198 474 -193
rect 552 -193 553 -189
rect 557 -193 558 -189
rect 594 -188 598 -159
rect 608 -162 612 -155
rect 608 -163 613 -162
rect 608 -167 609 -163
rect 616 -163 620 -142
rect 623 -148 636 -147
rect 623 -152 626 -148
rect 630 -152 632 -148
rect 623 -153 636 -152
rect 623 -160 629 -153
rect 639 -159 643 -142
rect 616 -167 619 -163
rect 623 -167 624 -163
rect 628 -167 629 -163
rect 633 -167 634 -163
rect 639 -164 643 -163
rect 608 -168 613 -167
rect 608 -176 612 -168
rect 628 -172 634 -167
rect 615 -176 616 -172
rect 620 -176 634 -172
rect 640 -173 644 -171
rect 565 -191 569 -190
rect 574 -192 575 -188
rect 579 -192 598 -188
rect 602 -179 612 -176
rect 602 -191 605 -179
rect 552 -198 558 -193
rect 608 -185 612 -179
rect 608 -186 613 -185
rect 608 -190 609 -186
rect 613 -190 620 -187
rect 608 -193 620 -190
rect 624 -189 628 -176
rect 640 -180 644 -177
rect 631 -184 635 -180
rect 639 -184 644 -180
rect 631 -185 644 -184
rect 624 -193 638 -189
rect 642 -193 643 -189
rect 375 -202 378 -198
rect 382 -202 388 -198
rect 392 -202 456 -198
rect 460 -202 509 -198
rect 513 -202 540 -198
rect 544 -202 593 -198
rect 597 -202 610 -198
rect 614 -202 620 -198
rect 624 -199 648 -198
rect 624 -202 640 -199
rect 375 -203 640 -202
rect 360 -205 640 -203
rect 646 -205 648 -199
rect 360 -206 648 -205
rect 360 -207 376 -206
rect 465 -208 509 -206
rect 465 -212 471 -208
rect 475 -212 499 -208
rect 503 -212 509 -208
rect 362 -231 430 -227
rect 171 -258 176 -257
rect 140 -264 141 -260
rect 145 -264 160 -260
rect 163 -262 171 -260
rect 175 -262 176 -258
rect 306 -259 333 -255
rect 163 -264 176 -262
rect 158 -270 159 -267
rect 136 -271 159 -270
rect 163 -270 164 -267
rect 163 -271 170 -270
rect 136 -274 170 -271
rect 174 -274 180 -270
rect 136 -275 180 -274
rect 341 -273 346 -253
rect 444 -254 447 -219
rect 469 -220 475 -212
rect 469 -224 470 -220
rect 474 -224 475 -220
rect 480 -220 484 -219
rect 489 -220 495 -212
rect 489 -224 490 -220
rect 494 -224 495 -220
rect 500 -220 505 -217
rect 545 -219 629 -216
rect 504 -224 505 -220
rect 480 -227 484 -224
rect 500 -225 505 -224
rect 480 -231 497 -227
rect 469 -243 473 -233
rect 477 -238 482 -234
rect 493 -235 497 -231
rect 477 -246 483 -242
rect 487 -246 490 -242
rect 477 -252 481 -246
rect 493 -250 497 -239
rect 464 -255 481 -252
rect 485 -254 497 -250
rect 501 -231 505 -225
rect 501 -234 652 -231
rect 656 -234 657 -231
rect 485 -258 489 -254
rect 501 -255 505 -234
rect 669 -250 673 -142
rect 703 -159 707 -152
rect 703 -160 708 -159
rect 703 -164 704 -160
rect 711 -160 715 -139
rect 718 -145 731 -144
rect 718 -149 721 -145
rect 725 -149 727 -145
rect 718 -150 731 -149
rect 718 -157 724 -150
rect 734 -156 738 -139
rect 804 -139 816 -138
rect 820 -138 900 -135
rect 820 -139 884 -138
rect 781 -150 793 -144
rect 800 -145 804 -142
rect 888 -139 900 -138
rect 904 -139 937 -135
rect 941 -139 951 -135
rect 955 -139 965 -135
rect 969 -139 975 -135
rect 814 -148 836 -144
rect 840 -148 841 -144
rect 854 -145 877 -144
rect 814 -149 818 -148
rect 854 -149 870 -145
rect 874 -149 877 -145
rect 800 -150 804 -149
rect 781 -153 786 -150
rect 781 -154 782 -153
rect 711 -164 714 -160
rect 718 -164 719 -160
rect 723 -164 724 -160
rect 728 -164 729 -160
rect 734 -161 738 -160
rect 703 -165 708 -164
rect 703 -173 707 -165
rect 723 -169 729 -164
rect 710 -173 711 -169
rect 715 -173 729 -169
rect 735 -171 739 -168
rect 703 -182 707 -177
rect 703 -183 708 -182
rect 703 -187 704 -183
rect 708 -187 715 -184
rect 703 -190 715 -187
rect 719 -186 723 -173
rect 735 -177 739 -175
rect 726 -181 730 -177
rect 734 -181 739 -177
rect 726 -182 739 -181
rect 748 -186 751 -167
rect 719 -190 733 -186
rect 737 -190 738 -186
rect 749 -190 751 -186
rect 762 -188 766 -159
rect 773 -157 782 -154
rect 807 -153 818 -149
rect 807 -157 811 -153
rect 825 -156 826 -152
rect 830 -156 841 -152
rect 773 -171 776 -157
rect 781 -158 786 -157
rect 790 -159 811 -157
rect 782 -163 790 -162
rect 794 -161 811 -159
rect 782 -166 794 -163
rect 782 -178 786 -166
rect 807 -168 811 -161
rect 815 -163 816 -159
rect 820 -160 821 -159
rect 820 -163 832 -160
rect 815 -164 832 -163
rect 828 -167 832 -164
rect 828 -168 833 -167
rect 796 -174 802 -169
rect 807 -172 819 -168
rect 823 -172 824 -168
rect 828 -172 829 -168
rect 796 -176 798 -174
rect 789 -178 798 -176
rect 828 -173 833 -172
rect 837 -172 841 -156
rect 828 -177 832 -173
rect 789 -182 802 -178
rect 808 -181 832 -177
rect 837 -176 839 -172
rect 782 -183 786 -182
rect 808 -183 812 -181
rect 762 -192 763 -188
rect 795 -190 796 -186
rect 800 -190 801 -186
rect 837 -185 841 -176
rect 808 -188 812 -187
rect 817 -189 818 -185
rect 822 -189 841 -185
rect 848 -188 851 -157
rect 795 -195 801 -190
rect 855 -195 859 -149
rect 865 -150 877 -149
rect 884 -145 888 -142
rect 898 -148 920 -144
rect 924 -148 925 -144
rect 898 -149 902 -148
rect 884 -150 888 -149
rect 865 -153 870 -150
rect 865 -157 866 -153
rect 891 -153 902 -149
rect 891 -157 895 -153
rect 909 -156 910 -152
rect 914 -156 925 -152
rect 865 -158 870 -157
rect 874 -159 895 -157
rect 866 -163 874 -162
rect 878 -161 895 -159
rect 866 -166 878 -163
rect 866 -178 870 -166
rect 891 -168 895 -161
rect 899 -163 900 -159
rect 904 -160 905 -159
rect 904 -163 916 -160
rect 899 -164 916 -163
rect 912 -167 916 -164
rect 912 -168 917 -167
rect 880 -174 886 -169
rect 891 -172 903 -168
rect 907 -172 908 -168
rect 912 -172 913 -168
rect 880 -176 882 -174
rect 873 -178 882 -176
rect 912 -173 917 -172
rect 912 -177 916 -173
rect 873 -182 886 -178
rect 892 -181 916 -177
rect 866 -183 870 -182
rect 892 -183 896 -181
rect 879 -190 880 -186
rect 884 -190 885 -186
rect 921 -185 925 -156
rect 935 -159 939 -152
rect 935 -160 940 -159
rect 935 -164 936 -160
rect 943 -160 947 -139
rect 950 -145 963 -144
rect 950 -149 953 -145
rect 957 -149 959 -145
rect 950 -150 963 -149
rect 950 -157 956 -150
rect 966 -156 970 -139
rect 943 -164 946 -160
rect 950 -164 951 -160
rect 955 -164 956 -160
rect 960 -164 961 -160
rect 966 -161 970 -160
rect 935 -165 940 -164
rect 935 -173 939 -165
rect 955 -169 961 -164
rect 942 -173 943 -169
rect 947 -173 961 -169
rect 967 -170 971 -168
rect 892 -188 896 -187
rect 901 -189 902 -185
rect 906 -189 925 -185
rect 929 -176 939 -173
rect 929 -188 932 -176
rect 879 -195 885 -190
rect 935 -182 939 -176
rect 935 -183 940 -182
rect 935 -187 936 -183
rect 940 -187 947 -184
rect 935 -190 947 -187
rect 951 -186 955 -173
rect 967 -177 971 -174
rect 958 -181 962 -177
rect 966 -181 971 -177
rect 958 -182 971 -181
rect 951 -190 965 -186
rect 969 -190 970 -186
rect 702 -196 705 -195
rect 700 -199 705 -196
rect 709 -199 715 -195
rect 719 -199 783 -195
rect 787 -199 836 -195
rect 840 -199 867 -195
rect 871 -199 920 -195
rect 924 -199 937 -195
rect 941 -199 947 -195
rect 951 -199 975 -195
rect 700 -201 975 -199
rect 687 -203 975 -201
rect 687 -204 704 -203
rect 687 -205 703 -204
rect 792 -205 836 -203
rect 792 -209 798 -205
rect 802 -209 826 -205
rect 830 -209 836 -205
rect 796 -217 802 -209
rect 500 -256 505 -255
rect 469 -262 470 -258
rect 474 -262 489 -258
rect 492 -260 500 -258
rect 504 -260 505 -256
rect 492 -262 505 -260
rect 630 -265 633 -251
rect 487 -268 488 -265
rect 465 -269 488 -268
rect 492 -268 493 -265
rect 630 -268 659 -265
rect 492 -269 499 -268
rect 465 -272 499 -269
rect 503 -272 509 -268
rect 465 -273 509 -272
rect 12 -278 180 -275
rect 12 -279 140 -278
rect 318 -279 333 -275
rect 137 -282 140 -279
rect 341 -276 509 -273
rect 341 -277 467 -276
rect 464 -280 467 -277
rect 12 -286 318 -282
rect 12 -290 48 -286
rect 52 -290 62 -286
rect 66 -290 76 -286
rect 80 -289 159 -286
rect 80 -290 143 -289
rect 12 -401 16 -290
rect 46 -310 50 -303
rect 46 -311 51 -310
rect 46 -315 47 -311
rect 54 -311 58 -290
rect 61 -296 74 -295
rect 61 -300 64 -296
rect 68 -300 70 -296
rect 61 -301 74 -300
rect 61 -308 67 -301
rect 77 -307 81 -290
rect 147 -290 159 -289
rect 163 -289 243 -286
rect 163 -290 227 -289
rect 124 -301 136 -295
rect 143 -296 147 -293
rect 231 -290 243 -289
rect 247 -290 280 -286
rect 284 -290 294 -286
rect 298 -290 308 -286
rect 312 -290 318 -286
rect 341 -284 647 -280
rect 341 -288 377 -284
rect 381 -288 391 -284
rect 395 -288 405 -284
rect 409 -287 488 -284
rect 409 -288 472 -287
rect 157 -299 179 -295
rect 183 -299 184 -295
rect 208 -296 220 -295
rect 196 -299 213 -296
rect 157 -300 161 -299
rect 143 -301 147 -300
rect 124 -304 129 -301
rect 124 -305 125 -304
rect 54 -315 57 -311
rect 61 -315 62 -311
rect 66 -315 67 -311
rect 71 -315 72 -311
rect 77 -312 81 -311
rect 116 -308 125 -305
rect 150 -304 161 -300
rect 150 -308 154 -304
rect 168 -307 169 -303
rect 173 -307 184 -303
rect 46 -316 51 -315
rect 46 -324 50 -316
rect 66 -320 72 -315
rect 53 -324 54 -320
rect 58 -324 72 -320
rect 78 -322 82 -319
rect 116 -322 119 -308
rect 124 -309 129 -308
rect 133 -310 154 -308
rect 46 -333 50 -328
rect 46 -334 51 -333
rect 46 -338 47 -334
rect 51 -338 58 -335
rect 46 -341 58 -338
rect 62 -337 66 -324
rect 125 -314 133 -313
rect 137 -312 154 -310
rect 125 -317 137 -314
rect 78 -328 82 -326
rect 69 -332 73 -328
rect 77 -332 82 -328
rect 69 -333 82 -332
rect 125 -329 129 -317
rect 150 -319 154 -312
rect 158 -314 159 -310
rect 163 -311 164 -310
rect 163 -314 175 -311
rect 158 -315 175 -314
rect 171 -318 175 -315
rect 171 -319 176 -318
rect 139 -325 145 -320
rect 150 -323 162 -319
rect 166 -323 167 -319
rect 171 -323 172 -319
rect 139 -327 141 -325
rect 132 -329 141 -327
rect 171 -324 176 -323
rect 180 -323 184 -307
rect 171 -328 175 -324
rect 132 -333 145 -329
rect 151 -332 175 -328
rect 180 -327 182 -323
rect 125 -334 129 -333
rect 151 -334 155 -332
rect 62 -341 76 -337
rect 80 -341 81 -337
rect 138 -341 139 -337
rect 143 -341 144 -337
rect 180 -336 184 -327
rect 151 -339 155 -338
rect 160 -340 161 -336
rect 165 -340 184 -336
rect 196 -339 199 -299
rect 208 -300 213 -299
rect 217 -300 220 -296
rect 208 -301 220 -300
rect 227 -296 231 -293
rect 241 -299 263 -295
rect 267 -299 268 -295
rect 241 -300 245 -299
rect 227 -301 231 -300
rect 208 -304 213 -301
rect 208 -308 209 -304
rect 234 -304 245 -300
rect 234 -308 238 -304
rect 252 -307 253 -303
rect 257 -307 268 -303
rect 208 -309 213 -308
rect 217 -310 238 -308
rect 264 -309 268 -307
rect 209 -314 217 -313
rect 221 -312 238 -310
rect 209 -317 221 -314
rect 209 -329 213 -317
rect 234 -319 238 -312
rect 242 -314 243 -310
rect 247 -311 248 -310
rect 247 -314 259 -311
rect 242 -315 259 -314
rect 255 -318 259 -315
rect 264 -312 271 -309
rect 278 -310 282 -303
rect 278 -311 283 -310
rect 255 -319 260 -318
rect 223 -325 229 -320
rect 234 -323 246 -319
rect 250 -323 251 -319
rect 255 -323 256 -319
rect 223 -327 225 -325
rect 216 -329 225 -327
rect 255 -324 260 -323
rect 255 -328 259 -324
rect 216 -333 229 -329
rect 235 -332 259 -328
rect 209 -334 213 -333
rect 235 -334 239 -332
rect 138 -346 144 -341
rect 222 -341 223 -337
rect 227 -341 228 -337
rect 264 -336 268 -312
rect 278 -315 279 -311
rect 286 -311 290 -290
rect 293 -296 306 -295
rect 293 -300 296 -296
rect 300 -300 302 -296
rect 293 -301 306 -300
rect 293 -308 299 -301
rect 309 -307 313 -290
rect 322 -308 333 -305
rect 286 -315 289 -311
rect 293 -315 294 -311
rect 298 -315 299 -311
rect 303 -315 304 -311
rect 309 -312 313 -311
rect 278 -316 283 -315
rect 278 -324 282 -316
rect 298 -320 304 -315
rect 285 -324 286 -320
rect 290 -324 304 -320
rect 310 -321 314 -319
rect 235 -339 239 -338
rect 244 -340 245 -336
rect 249 -340 268 -336
rect 272 -327 282 -324
rect 272 -339 275 -327
rect 222 -346 228 -341
rect 278 -333 282 -327
rect 278 -334 283 -333
rect 278 -338 279 -334
rect 283 -338 290 -335
rect 278 -341 290 -338
rect 294 -337 298 -324
rect 310 -328 314 -325
rect 301 -332 305 -328
rect 309 -332 314 -328
rect 301 -333 314 -332
rect 294 -341 308 -337
rect 312 -341 313 -337
rect 45 -350 48 -346
rect 52 -350 58 -346
rect 62 -350 126 -346
rect 130 -350 179 -346
rect 183 -350 210 -346
rect 214 -350 263 -346
rect 267 -350 280 -346
rect 284 -350 290 -346
rect 294 -350 313 -346
rect 45 -353 313 -350
rect 45 -354 318 -353
rect 135 -356 179 -354
rect 135 -360 141 -356
rect 145 -360 169 -356
rect 173 -360 179 -356
rect 139 -368 145 -360
rect 139 -372 140 -368
rect 144 -372 145 -368
rect 150 -368 154 -367
rect 159 -368 165 -360
rect 266 -363 307 -360
rect 159 -372 160 -368
rect 164 -372 165 -368
rect 170 -368 175 -365
rect 174 -372 175 -368
rect 150 -375 154 -372
rect 170 -373 175 -372
rect 150 -379 167 -375
rect 139 -391 143 -381
rect 147 -386 152 -382
rect 163 -383 167 -379
rect 147 -394 153 -390
rect 157 -394 160 -390
rect 11 -421 16 -401
rect 147 -400 151 -394
rect 163 -398 167 -387
rect 134 -403 151 -400
rect 155 -402 167 -398
rect 171 -385 175 -373
rect 263 -381 286 -378
rect 291 -381 292 -378
rect 171 -388 250 -385
rect 155 -406 159 -402
rect 171 -403 175 -388
rect 170 -404 175 -403
rect 139 -410 140 -406
rect 144 -410 159 -406
rect 162 -408 170 -406
rect 174 -408 175 -404
rect 247 -403 250 -388
rect 247 -406 293 -403
rect 162 -410 175 -408
rect 157 -416 158 -413
rect 135 -417 158 -416
rect 162 -416 163 -413
rect 162 -417 169 -416
rect 135 -420 169 -417
rect 173 -420 179 -416
rect 135 -421 179 -420
rect 11 -424 179 -421
rect 11 -425 135 -424
rect 304 -464 307 -363
rect 316 -382 332 -378
rect 341 -399 345 -288
rect 375 -308 379 -301
rect 375 -309 380 -308
rect 375 -313 376 -309
rect 383 -309 387 -288
rect 390 -294 403 -293
rect 390 -298 393 -294
rect 397 -298 399 -294
rect 390 -299 403 -298
rect 390 -306 396 -299
rect 406 -305 410 -288
rect 476 -288 488 -287
rect 492 -287 572 -284
rect 492 -288 556 -287
rect 453 -299 465 -293
rect 472 -294 476 -291
rect 560 -288 572 -287
rect 576 -288 609 -284
rect 613 -288 623 -284
rect 627 -288 637 -284
rect 641 -288 647 -284
rect 486 -297 508 -293
rect 512 -297 513 -293
rect 537 -294 549 -293
rect 486 -298 490 -297
rect 472 -299 476 -298
rect 453 -302 458 -299
rect 453 -303 454 -302
rect 383 -313 386 -309
rect 390 -313 391 -309
rect 395 -313 396 -309
rect 400 -313 401 -309
rect 406 -310 410 -309
rect 445 -306 454 -303
rect 479 -302 490 -298
rect 537 -298 542 -294
rect 546 -298 549 -294
rect 537 -299 549 -298
rect 556 -294 560 -291
rect 570 -297 592 -293
rect 596 -297 597 -293
rect 570 -298 574 -297
rect 556 -299 560 -298
rect 479 -306 483 -302
rect 497 -305 498 -301
rect 502 -305 513 -301
rect 375 -314 380 -313
rect 375 -322 379 -314
rect 395 -318 401 -313
rect 382 -322 383 -318
rect 387 -322 401 -318
rect 407 -320 411 -317
rect 375 -331 379 -326
rect 375 -332 380 -331
rect 375 -336 376 -332
rect 380 -336 387 -333
rect 375 -339 387 -336
rect 391 -335 395 -322
rect 407 -326 411 -324
rect 398 -330 402 -326
rect 406 -330 411 -326
rect 398 -331 411 -330
rect 391 -339 405 -335
rect 409 -339 410 -335
rect 435 -337 438 -317
rect 445 -320 448 -306
rect 453 -307 458 -306
rect 462 -308 483 -306
rect 454 -312 462 -311
rect 466 -310 483 -308
rect 454 -315 466 -312
rect 454 -327 458 -315
rect 479 -317 483 -310
rect 487 -312 488 -308
rect 492 -309 493 -308
rect 492 -312 504 -309
rect 487 -313 504 -312
rect 500 -316 504 -313
rect 500 -317 505 -316
rect 468 -323 474 -318
rect 479 -321 491 -317
rect 495 -321 496 -317
rect 500 -321 501 -317
rect 468 -325 470 -323
rect 461 -327 470 -325
rect 500 -322 505 -321
rect 509 -321 513 -305
rect 537 -302 542 -299
rect 537 -306 538 -302
rect 563 -302 574 -298
rect 563 -306 567 -302
rect 581 -305 582 -301
rect 586 -305 597 -301
rect 537 -307 542 -306
rect 546 -308 567 -306
rect 538 -312 546 -311
rect 550 -310 567 -308
rect 538 -315 550 -312
rect 500 -326 504 -322
rect 461 -331 474 -327
rect 480 -330 504 -326
rect 509 -325 511 -321
rect 454 -332 458 -331
rect 480 -332 484 -330
rect 467 -339 468 -335
rect 472 -339 473 -335
rect 509 -334 513 -325
rect 538 -327 542 -315
rect 563 -317 567 -310
rect 571 -312 572 -308
rect 576 -309 577 -308
rect 576 -312 588 -309
rect 571 -313 588 -312
rect 584 -316 588 -313
rect 593 -311 597 -305
rect 607 -308 611 -301
rect 607 -309 612 -308
rect 593 -314 600 -311
rect 607 -313 608 -309
rect 615 -309 619 -288
rect 622 -294 635 -293
rect 622 -298 625 -294
rect 629 -298 631 -294
rect 622 -299 635 -298
rect 622 -306 628 -299
rect 638 -305 642 -288
rect 615 -313 618 -309
rect 622 -313 623 -309
rect 627 -313 628 -309
rect 632 -313 633 -309
rect 638 -310 642 -309
rect 607 -314 612 -313
rect 584 -317 589 -316
rect 552 -323 558 -318
rect 563 -321 575 -317
rect 579 -321 580 -317
rect 584 -321 585 -317
rect 552 -325 554 -323
rect 545 -327 554 -325
rect 584 -322 589 -321
rect 584 -326 588 -322
rect 545 -331 558 -327
rect 564 -330 588 -326
rect 538 -332 542 -331
rect 564 -332 568 -330
rect 480 -337 484 -336
rect 489 -338 490 -334
rect 494 -338 513 -334
rect 467 -344 473 -339
rect 551 -339 552 -335
rect 556 -339 557 -335
rect 593 -334 597 -314
rect 607 -322 611 -314
rect 627 -318 633 -313
rect 614 -322 615 -318
rect 619 -322 633 -318
rect 639 -319 643 -317
rect 564 -337 568 -336
rect 573 -338 574 -334
rect 578 -338 597 -334
rect 601 -325 611 -322
rect 601 -337 604 -325
rect 551 -344 557 -339
rect 607 -331 611 -325
rect 607 -332 612 -331
rect 607 -336 608 -332
rect 612 -336 619 -333
rect 607 -339 619 -336
rect 623 -335 627 -322
rect 639 -326 643 -323
rect 630 -330 634 -326
rect 638 -330 643 -326
rect 630 -331 643 -330
rect 623 -339 637 -335
rect 641 -339 642 -335
rect 374 -348 377 -344
rect 381 -348 387 -344
rect 391 -348 455 -344
rect 459 -348 508 -344
rect 512 -348 539 -344
rect 543 -348 592 -344
rect 596 -348 609 -344
rect 613 -348 619 -344
rect 623 -348 647 -344
rect 355 -351 640 -348
rect 374 -352 640 -351
rect 644 -352 647 -348
rect 464 -354 508 -352
rect 384 -356 446 -355
rect 388 -358 446 -356
rect 388 -359 424 -358
rect 464 -358 470 -354
rect 474 -358 498 -354
rect 502 -358 508 -354
rect 435 -363 438 -361
rect 468 -366 474 -358
rect 363 -374 411 -371
rect 435 -381 438 -367
rect 468 -370 469 -366
rect 473 -370 474 -366
rect 479 -366 483 -365
rect 488 -366 494 -358
rect 634 -356 638 -355
rect 592 -359 638 -356
rect 488 -370 489 -366
rect 493 -370 494 -366
rect 499 -366 504 -363
rect 503 -370 504 -366
rect 479 -373 483 -370
rect 499 -371 504 -370
rect 479 -377 496 -373
rect 317 -406 332 -403
rect 340 -419 345 -399
rect 385 -411 389 -383
rect 407 -385 435 -382
rect 407 -411 411 -385
rect 468 -389 472 -379
rect 476 -384 481 -380
rect 492 -381 496 -377
rect 476 -392 482 -388
rect 486 -392 489 -388
rect 476 -398 480 -392
rect 492 -396 496 -385
rect 463 -401 480 -398
rect 484 -400 496 -396
rect 484 -404 488 -400
rect 500 -401 504 -371
rect 531 -375 613 -370
rect 634 -390 638 -359
rect 637 -393 638 -390
rect 499 -402 504 -401
rect 468 -408 469 -404
rect 473 -408 488 -404
rect 491 -406 499 -404
rect 503 -404 504 -402
rect 503 -406 508 -404
rect 491 -408 508 -406
rect 486 -414 487 -411
rect 464 -415 487 -414
rect 491 -414 492 -411
rect 491 -415 498 -414
rect 464 -418 498 -415
rect 502 -418 508 -414
rect 464 -419 508 -418
rect 340 -422 508 -419
rect 340 -423 464 -422
rect 453 -430 457 -423
rect 336 -432 380 -430
rect 429 -432 473 -430
rect 516 -432 560 -430
rect 336 -434 560 -432
rect 336 -438 342 -434
rect 346 -435 435 -434
rect 346 -438 380 -435
rect 429 -438 435 -435
rect 439 -435 522 -434
rect 439 -438 473 -435
rect 516 -438 522 -435
rect 526 -438 560 -434
rect 656 -438 659 -268
rect 668 -270 673 -250
rect 677 -222 680 -221
rect 677 -225 712 -222
rect 796 -221 797 -217
rect 801 -221 802 -217
rect 807 -217 811 -216
rect 816 -217 822 -209
rect 816 -221 817 -217
rect 821 -221 822 -217
rect 827 -217 832 -214
rect 831 -221 832 -217
rect 677 -262 680 -225
rect 688 -234 755 -231
rect 759 -234 760 -231
rect 765 -262 769 -222
rect 807 -224 811 -221
rect 827 -222 832 -221
rect 807 -228 824 -224
rect 777 -256 780 -229
rect 796 -240 800 -230
rect 804 -235 809 -231
rect 820 -232 824 -228
rect 804 -243 810 -239
rect 814 -243 817 -239
rect 804 -249 808 -243
rect 820 -247 824 -236
rect 791 -252 808 -249
rect 812 -251 824 -247
rect 828 -226 832 -222
rect 828 -229 840 -226
rect 812 -255 816 -251
rect 828 -252 832 -229
rect 848 -250 851 -235
rect 827 -253 832 -252
rect 796 -259 797 -255
rect 801 -259 816 -255
rect 819 -257 827 -255
rect 831 -257 832 -253
rect 819 -259 832 -257
rect 677 -263 686 -262
rect 677 -267 696 -263
rect 700 -267 705 -263
rect 814 -265 815 -262
rect 765 -267 769 -266
rect 792 -266 815 -265
rect 819 -265 820 -262
rect 847 -263 852 -250
rect 819 -266 826 -265
rect 792 -269 826 -266
rect 830 -269 836 -265
rect 792 -270 836 -269
rect 997 -267 1001 -266
rect 668 -273 836 -270
rect 964 -270 1002 -267
rect 1012 -270 1015 -129
rect 1192 -131 1197 -128
rect 1298 -131 1302 -128
rect 1124 -134 1373 -131
rect 1124 -139 1127 -134
rect 1170 -140 1173 -134
rect 1224 -140 1227 -134
rect 1280 -140 1283 -134
rect 1334 -140 1337 -134
rect 1021 -186 1025 -147
rect 1158 -151 1161 -143
rect 1158 -155 1159 -151
rect 1141 -164 1144 -161
rect 1158 -177 1161 -155
rect 1204 -157 1207 -144
rect 1204 -160 1214 -157
rect 1246 -160 1249 -156
rect 1258 -154 1261 -144
rect 1258 -157 1277 -154
rect 1306 -154 1309 -153
rect 1173 -164 1175 -161
rect 1195 -164 1196 -161
rect 1204 -169 1207 -160
rect 1171 -172 1207 -169
rect 1171 -177 1174 -172
rect 1204 -177 1207 -172
rect 1211 -169 1214 -160
rect 1225 -164 1229 -162
rect 1246 -163 1250 -160
rect 1225 -165 1232 -164
rect 1258 -169 1261 -157
rect 1308 -158 1309 -154
rect 1306 -160 1309 -158
rect 1282 -164 1285 -161
rect 1314 -164 1317 -144
rect 1340 -151 1341 -147
rect 1338 -160 1341 -151
rect 1368 -155 1371 -144
rect 1338 -163 1339 -160
rect 1357 -164 1360 -162
rect 1357 -165 1363 -164
rect 1314 -169 1317 -168
rect 1368 -169 1371 -159
rect 1225 -172 1261 -169
rect 1225 -177 1228 -172
rect 1258 -177 1261 -172
rect 1281 -172 1317 -169
rect 1281 -177 1284 -172
rect 1314 -177 1317 -172
rect 1335 -172 1371 -169
rect 1335 -177 1338 -172
rect 1368 -177 1371 -172
rect 1124 -200 1127 -181
rect 1187 -200 1190 -181
rect 1197 -200 1200 -195
rect 1241 -200 1244 -181
rect 1251 -200 1254 -195
rect 1297 -200 1300 -181
rect 1307 -200 1310 -195
rect 1351 -200 1354 -181
rect 1361 -200 1364 -195
rect 1382 -200 1387 -59
rect 1407 -141 1412 -38
rect 1122 -201 1387 -200
rect 1019 -203 1387 -201
rect 1019 -204 1385 -203
rect 1035 -223 1038 -204
rect 1080 -221 1084 -219
rect 1118 -223 1121 -204
rect 1132 -212 1161 -209
rect 1080 -238 1084 -227
rect 1063 -242 1066 -239
rect 1080 -248 1083 -238
rect 1135 -243 1138 -240
rect 1080 -252 1081 -248
rect 1152 -249 1155 -227
rect 1158 -239 1161 -212
rect 1181 -223 1184 -204
rect 1191 -209 1194 -204
rect 1235 -223 1238 -204
rect 1245 -209 1248 -204
rect 1291 -223 1294 -204
rect 1301 -209 1304 -204
rect 1345 -223 1348 -204
rect 1355 -209 1358 -204
rect 1165 -232 1168 -227
rect 1198 -232 1201 -227
rect 1165 -235 1201 -232
rect 1158 -242 1163 -239
rect 1167 -243 1169 -240
rect 1189 -243 1190 -240
rect 1198 -244 1201 -235
rect 1219 -232 1222 -227
rect 1252 -232 1255 -227
rect 1219 -235 1255 -232
rect 1275 -232 1278 -227
rect 1308 -232 1311 -227
rect 1275 -235 1311 -232
rect 1329 -232 1332 -227
rect 1362 -232 1365 -227
rect 1329 -235 1365 -232
rect 1205 -244 1208 -235
rect 1219 -240 1226 -239
rect 1219 -242 1223 -240
rect 1240 -244 1244 -241
rect 1198 -247 1208 -244
rect 1080 -260 1083 -252
rect 1152 -253 1153 -249
rect 1152 -261 1155 -253
rect 1198 -260 1201 -247
rect 1240 -248 1243 -244
rect 1252 -247 1255 -235
rect 1308 -236 1311 -235
rect 1276 -243 1279 -240
rect 1252 -250 1271 -247
rect 1252 -260 1255 -250
rect 1300 -246 1303 -244
rect 1288 -254 1291 -248
rect 1302 -250 1303 -246
rect 1300 -251 1303 -250
rect 1265 -257 1291 -254
rect 1308 -260 1311 -240
rect 1332 -244 1333 -241
rect 1351 -240 1357 -239
rect 1351 -242 1354 -240
rect 1332 -253 1335 -244
rect 1362 -245 1365 -235
rect 1334 -257 1335 -253
rect 1362 -260 1365 -249
rect 1046 -270 1049 -264
rect 1118 -270 1121 -265
rect 1164 -270 1167 -264
rect 1218 -270 1221 -264
rect 1274 -270 1277 -264
rect 1328 -270 1331 -264
rect 668 -274 792 -273
rect 797 -277 800 -273
rect 668 -281 974 -277
rect 668 -285 704 -281
rect 708 -285 718 -281
rect 722 -285 732 -281
rect 736 -284 815 -281
rect 736 -285 799 -284
rect 668 -396 672 -285
rect 702 -305 706 -298
rect 702 -306 707 -305
rect 702 -310 703 -306
rect 710 -306 714 -285
rect 717 -291 730 -290
rect 717 -295 720 -291
rect 724 -295 726 -291
rect 717 -296 730 -295
rect 717 -303 723 -296
rect 733 -302 737 -285
rect 803 -285 815 -284
rect 819 -284 899 -281
rect 819 -285 883 -284
rect 780 -296 792 -290
rect 799 -291 803 -288
rect 887 -285 899 -284
rect 903 -285 936 -281
rect 940 -285 950 -281
rect 954 -285 964 -281
rect 968 -285 974 -281
rect 813 -294 835 -290
rect 839 -294 840 -290
rect 864 -291 876 -290
rect 813 -295 817 -294
rect 799 -296 803 -295
rect 780 -299 785 -296
rect 710 -310 713 -306
rect 717 -310 718 -306
rect 722 -310 723 -306
rect 727 -310 728 -306
rect 733 -307 737 -306
rect 780 -300 781 -299
rect 702 -311 707 -310
rect 702 -319 706 -311
rect 722 -315 728 -310
rect 709 -319 710 -315
rect 714 -319 728 -315
rect 734 -317 738 -314
rect 702 -328 706 -323
rect 702 -329 707 -328
rect 702 -333 703 -329
rect 707 -333 714 -330
rect 702 -336 714 -333
rect 718 -332 722 -319
rect 734 -323 738 -321
rect 725 -327 729 -323
rect 733 -327 738 -323
rect 725 -328 738 -327
rect 751 -329 755 -304
rect 772 -303 781 -300
rect 806 -299 817 -295
rect 864 -295 869 -291
rect 873 -295 876 -291
rect 864 -296 876 -295
rect 883 -291 887 -288
rect 897 -294 919 -290
rect 923 -294 924 -290
rect 897 -295 901 -294
rect 883 -296 887 -295
rect 806 -303 810 -299
rect 824 -302 825 -298
rect 829 -302 840 -298
rect 772 -317 775 -303
rect 780 -304 785 -303
rect 789 -305 810 -303
rect 781 -309 789 -308
rect 793 -307 810 -305
rect 781 -312 793 -309
rect 781 -324 785 -312
rect 806 -314 810 -307
rect 814 -309 815 -305
rect 819 -306 820 -305
rect 819 -309 831 -306
rect 814 -310 831 -309
rect 827 -313 831 -310
rect 827 -314 832 -313
rect 795 -320 801 -315
rect 806 -318 818 -314
rect 822 -318 823 -314
rect 827 -318 828 -314
rect 795 -322 797 -320
rect 781 -329 785 -328
rect 788 -324 797 -322
rect 827 -319 832 -318
rect 836 -318 840 -302
rect 864 -299 869 -296
rect 864 -303 865 -299
rect 890 -299 901 -295
rect 890 -303 894 -299
rect 908 -302 909 -298
rect 913 -302 924 -298
rect 864 -304 869 -303
rect 873 -305 894 -303
rect 865 -309 873 -308
rect 877 -307 894 -305
rect 865 -312 877 -309
rect 827 -323 831 -319
rect 788 -328 801 -324
rect 807 -327 831 -323
rect 836 -322 838 -318
rect 718 -336 732 -332
rect 736 -336 737 -332
rect 753 -332 755 -329
rect 788 -333 791 -328
rect 807 -329 811 -327
rect 777 -337 791 -333
rect 794 -336 795 -332
rect 799 -336 800 -332
rect 836 -331 840 -322
rect 865 -324 869 -312
rect 890 -314 894 -307
rect 898 -309 899 -305
rect 903 -306 904 -305
rect 903 -309 915 -306
rect 898 -310 915 -309
rect 911 -313 915 -310
rect 920 -307 924 -302
rect 934 -305 938 -298
rect 934 -306 939 -305
rect 920 -311 927 -307
rect 934 -310 935 -306
rect 942 -306 946 -285
rect 949 -291 962 -290
rect 949 -295 952 -291
rect 956 -295 958 -291
rect 949 -296 962 -295
rect 949 -303 955 -296
rect 965 -302 969 -285
rect 942 -310 945 -306
rect 949 -310 950 -306
rect 954 -310 955 -306
rect 959 -310 960 -306
rect 965 -307 969 -306
rect 934 -311 939 -310
rect 911 -314 916 -313
rect 879 -320 885 -315
rect 890 -318 902 -314
rect 906 -318 907 -314
rect 911 -318 912 -314
rect 879 -322 881 -320
rect 872 -324 881 -322
rect 911 -319 916 -318
rect 911 -323 915 -319
rect 872 -328 885 -324
rect 891 -327 915 -323
rect 865 -329 869 -328
rect 891 -329 895 -327
rect 807 -334 811 -333
rect 816 -335 817 -331
rect 821 -335 840 -331
rect 777 -341 781 -337
rect 794 -341 800 -336
rect 878 -336 879 -332
rect 883 -336 884 -332
rect 920 -331 924 -311
rect 934 -319 938 -311
rect 954 -315 960 -310
rect 941 -319 942 -315
rect 946 -319 960 -315
rect 966 -316 970 -314
rect 891 -334 895 -333
rect 900 -335 901 -331
rect 905 -335 924 -331
rect 928 -322 938 -319
rect 928 -334 931 -322
rect 878 -341 884 -336
rect 934 -328 938 -322
rect 934 -329 939 -328
rect 934 -333 935 -329
rect 939 -333 946 -330
rect 934 -336 946 -333
rect 950 -332 954 -319
rect 966 -323 970 -320
rect 957 -327 961 -323
rect 965 -327 970 -323
rect 957 -328 970 -327
rect 950 -336 964 -332
rect 968 -336 969 -332
rect 701 -344 704 -341
rect 700 -345 704 -344
rect 708 -345 714 -341
rect 718 -345 782 -341
rect 786 -345 835 -341
rect 839 -345 866 -341
rect 870 -345 919 -341
rect 923 -345 936 -341
rect 940 -345 946 -341
rect 950 -345 974 -341
rect 700 -347 974 -345
rect 681 -348 974 -347
rect 684 -349 974 -348
rect 684 -350 703 -349
rect 791 -351 835 -349
rect 791 -355 797 -351
rect 801 -355 825 -351
rect 829 -355 835 -351
rect 738 -357 742 -356
rect 682 -375 711 -370
rect 667 -416 672 -396
rect 738 -398 742 -361
rect 795 -363 801 -355
rect 795 -367 796 -363
rect 800 -367 801 -363
rect 806 -363 810 -362
rect 815 -363 821 -355
rect 815 -367 816 -363
rect 820 -367 821 -363
rect 826 -363 831 -360
rect 830 -367 831 -363
rect 806 -370 810 -367
rect 826 -368 831 -367
rect 806 -374 823 -370
rect 754 -402 757 -383
rect 795 -386 799 -376
rect 803 -381 808 -377
rect 819 -378 823 -374
rect 827 -373 843 -368
rect 827 -378 831 -373
rect 803 -389 809 -385
rect 813 -389 816 -385
rect 803 -395 807 -389
rect 819 -393 823 -382
rect 826 -383 840 -378
rect 790 -398 807 -395
rect 811 -397 823 -393
rect 811 -401 815 -397
rect 827 -398 831 -383
rect 826 -399 831 -398
rect 795 -405 796 -401
rect 800 -405 815 -401
rect 818 -403 826 -401
rect 830 -403 831 -399
rect 818 -405 831 -403
rect 911 -408 915 -401
rect 813 -411 814 -408
rect 791 -412 814 -411
rect 818 -411 819 -408
rect 818 -412 825 -411
rect 791 -415 825 -412
rect 829 -415 835 -411
rect 791 -416 835 -415
rect 907 -416 916 -408
rect 667 -419 835 -416
rect 997 -418 1001 -270
rect 1011 -273 1364 -270
rect 1012 -412 1015 -273
rect 1190 -276 1195 -273
rect 1296 -276 1300 -273
rect 1122 -279 1368 -276
rect 1122 -284 1125 -279
rect 1168 -285 1171 -279
rect 1222 -285 1225 -279
rect 1278 -285 1281 -279
rect 1156 -296 1159 -288
rect 1156 -300 1157 -296
rect 1139 -309 1142 -306
rect 1156 -322 1159 -300
rect 1202 -302 1205 -289
rect 1202 -305 1212 -302
rect 1244 -305 1247 -301
rect 1256 -299 1259 -289
rect 1256 -302 1275 -299
rect 1304 -299 1307 -298
rect 1171 -309 1173 -306
rect 1193 -309 1194 -306
rect 1202 -314 1205 -305
rect 1169 -317 1205 -314
rect 1169 -322 1172 -317
rect 1202 -322 1205 -317
rect 1209 -314 1212 -305
rect 1223 -309 1227 -307
rect 1244 -308 1248 -305
rect 1223 -310 1230 -309
rect 1256 -314 1259 -302
rect 1306 -303 1307 -299
rect 1304 -305 1307 -303
rect 1280 -309 1283 -306
rect 1312 -309 1315 -289
rect 1312 -314 1315 -313
rect 1223 -317 1259 -314
rect 1223 -322 1226 -317
rect 1256 -322 1259 -317
rect 1279 -317 1315 -314
rect 1279 -322 1282 -317
rect 1312 -322 1315 -317
rect 1122 -343 1125 -326
rect 1185 -343 1188 -326
rect 1195 -343 1198 -340
rect 1239 -343 1242 -326
rect 1249 -343 1252 -340
rect 1295 -343 1298 -326
rect 1323 -335 1326 -286
rect 1332 -285 1335 -279
rect 1338 -296 1339 -292
rect 1336 -305 1339 -296
rect 1366 -300 1369 -289
rect 1336 -308 1337 -305
rect 1355 -309 1358 -307
rect 1355 -310 1361 -309
rect 1366 -314 1369 -304
rect 1333 -317 1369 -314
rect 1333 -322 1336 -317
rect 1366 -322 1369 -317
rect 1380 -301 1385 -204
rect 1435 -218 1441 19
rect 1498 -4 1502 115
rect 1633 113 1657 115
rect 1633 112 1674 113
rect 1521 109 1555 112
rect 1521 102 1525 109
rect 1538 79 1541 101
rect 1552 64 1555 109
rect 1633 108 1653 112
rect 1657 109 1674 112
rect 1678 109 1679 113
rect 1686 110 1688 114
rect 1692 110 1700 114
rect 1695 109 1700 110
rect 1633 98 1657 108
rect 1633 94 1653 98
rect 1633 90 1657 94
rect 1662 102 1663 106
rect 1667 102 1668 106
rect 1699 105 1700 109
rect 1662 100 1668 102
rect 1662 96 1663 100
rect 1667 99 1668 100
rect 1678 103 1691 104
rect 1682 99 1691 103
rect 1695 101 1700 105
rect 1704 112 1708 113
rect 1667 96 1675 99
rect 1678 98 1691 99
rect 1704 98 1708 108
rect 1662 93 1675 96
rect 1687 94 1708 98
rect 1713 94 1721 118
rect 1678 93 1682 94
rect 1633 89 1678 90
rect 1633 86 1682 89
rect 1687 90 1691 94
rect 1717 90 1721 94
rect 1569 83 1577 86
rect 1569 79 1573 83
rect 1569 73 1577 79
rect 1582 84 1595 85
rect 1582 80 1585 84
rect 1589 81 1595 84
rect 1599 84 1620 85
rect 1599 81 1608 84
rect 1589 80 1590 81
rect 1607 80 1608 81
rect 1612 81 1620 84
rect 1633 84 1657 86
rect 1687 85 1691 86
rect 1633 83 1653 84
rect 1612 80 1613 81
rect 1582 73 1588 80
rect 1637 80 1653 83
rect 1702 83 1708 90
rect 1677 82 1678 83
rect 1637 79 1657 80
rect 1599 77 1603 78
rect 1633 77 1657 79
rect 1670 79 1678 82
rect 1682 82 1683 83
rect 1700 82 1701 83
rect 1682 79 1701 82
rect 1705 79 1708 83
rect 1670 78 1708 79
rect 1713 84 1721 90
rect 1717 80 1721 84
rect 1569 69 1573 73
rect 1599 69 1603 73
rect 1608 74 1657 77
rect 1691 75 1694 78
rect 1612 73 1657 74
rect 1608 69 1612 70
rect 1569 5 1577 69
rect 1582 65 1603 69
rect 1615 67 1628 70
rect 1582 55 1586 65
rect 1599 64 1612 65
rect 1615 64 1623 67
rect 1582 50 1586 51
rect 1590 58 1595 62
rect 1599 60 1608 64
rect 1599 59 1612 60
rect 1622 63 1623 64
rect 1627 63 1628 67
rect 1622 61 1628 63
rect 1590 54 1591 58
rect 1622 57 1623 61
rect 1627 57 1628 61
rect 1633 69 1657 73
rect 1691 72 1706 75
rect 1637 65 1657 69
rect 1679 68 1682 71
rect 1633 55 1657 65
rect 1590 53 1595 54
rect 1590 49 1597 53
rect 1601 49 1604 53
rect 1611 50 1612 54
rect 1616 51 1633 54
rect 1637 51 1657 55
rect 1616 50 1657 51
rect 1633 47 1657 50
rect 1633 43 1653 47
rect 1585 40 1606 43
rect 1633 31 1657 43
rect 1662 67 1666 68
rect 1662 45 1666 63
rect 1670 64 1707 68
rect 1670 57 1674 64
rect 1685 59 1686 60
rect 1670 52 1674 53
rect 1678 56 1686 59
rect 1690 59 1691 60
rect 1690 56 1699 59
rect 1678 55 1699 56
rect 1678 48 1682 55
rect 1677 47 1682 48
rect 1662 41 1671 45
rect 1681 43 1682 47
rect 1677 42 1682 43
rect 1686 50 1690 51
rect 1667 38 1671 41
rect 1686 38 1690 46
rect 1667 34 1690 38
rect 1695 39 1699 55
rect 1703 49 1707 64
rect 1703 44 1707 45
rect 1713 67 1721 80
rect 1717 63 1721 67
rect 1695 35 1701 39
rect 1705 35 1706 39
rect 1588 28 1609 31
rect 1633 27 1656 31
rect 1660 27 1663 31
rect 1667 27 1668 31
rect 1601 12 1618 15
rect 1615 7 1618 12
rect 1614 6 1628 7
rect 1569 1 1573 5
rect 1589 2 1590 6
rect 1594 2 1610 6
rect 1614 2 1615 6
rect 1619 2 1628 6
rect 1499 -26 1507 -4
rect 1513 -9 1517 -8
rect 1513 -24 1517 -13
rect 1520 -16 1523 -3
rect 1569 -4 1577 1
rect 1563 -7 1577 -4
rect 1563 -8 1586 -7
rect 1532 -12 1542 -8
rect 1551 -9 1582 -8
rect 1555 -10 1582 -9
rect 1555 -13 1563 -10
rect 1551 -14 1563 -13
rect 1567 -12 1582 -10
rect 1567 -13 1586 -12
rect 1590 -8 1596 -1
rect 1606 -2 1610 2
rect 1606 -6 1609 -2
rect 1613 -6 1615 -2
rect 1622 -5 1628 2
rect 1590 -10 1603 -8
rect 1567 -14 1577 -13
rect 1590 -14 1594 -10
rect 1598 -14 1603 -10
rect 1520 -20 1533 -16
rect 1529 -22 1533 -20
rect 1537 -21 1541 -16
rect 1499 -27 1510 -26
rect 1499 -31 1506 -27
rect 1513 -28 1525 -24
rect 1499 -32 1510 -31
rect 1499 -38 1507 -32
rect 1499 -42 1503 -38
rect 1499 -48 1507 -42
rect 1513 -39 1517 -31
rect 1521 -32 1525 -28
rect 1544 -23 1551 -19
rect 1555 -23 1556 -19
rect 1529 -29 1533 -26
rect 1544 -32 1548 -23
rect 1563 -28 1577 -14
rect 1611 -19 1615 -6
rect 1633 -12 1657 27
rect 1675 21 1679 34
rect 1687 25 1692 29
rect 1696 25 1700 29
rect 1713 28 1721 63
rect 1687 23 1700 25
rect 1662 17 1668 20
rect 1675 17 1677 21
rect 1681 17 1684 21
rect 1662 13 1663 17
rect 1667 13 1668 17
rect 1680 13 1684 17
rect 1694 16 1700 23
rect 1704 27 1721 28
rect 1708 23 1721 27
rect 1704 22 1721 23
rect 1713 14 1721 22
rect 1662 9 1671 13
rect 1675 9 1676 13
rect 1680 9 1696 13
rect 1700 9 1701 13
rect 1717 10 1721 14
rect 1662 8 1676 9
rect 1666 -6 1705 -3
rect 1709 -6 1710 -3
rect 1622 -16 1623 -12
rect 1627 -16 1630 -12
rect 1634 -16 1657 -12
rect 1584 -24 1585 -20
rect 1589 -24 1595 -20
rect 1521 -36 1536 -32
rect 1540 -36 1548 -32
rect 1551 -29 1577 -28
rect 1555 -33 1577 -29
rect 1551 -34 1577 -33
rect 1563 -38 1577 -34
rect 1513 -43 1515 -39
rect 1519 -40 1520 -39
rect 1550 -40 1551 -39
rect 1519 -43 1537 -40
rect 1513 -44 1537 -43
rect 1541 -43 1551 -40
rect 1555 -43 1558 -39
rect 1541 -44 1558 -43
rect 1567 -42 1577 -38
rect 1563 -48 1577 -42
rect 1569 -52 1573 -48
rect 1569 -79 1577 -52
rect 1583 -30 1587 -29
rect 1583 -49 1587 -34
rect 1591 -40 1595 -24
rect 1600 -23 1623 -19
rect 1600 -31 1604 -23
rect 1619 -26 1623 -23
rect 1600 -36 1604 -35
rect 1608 -28 1613 -27
rect 1608 -32 1609 -28
rect 1619 -30 1628 -26
rect 1608 -33 1613 -32
rect 1608 -40 1612 -33
rect 1591 -41 1612 -40
rect 1591 -44 1600 -41
rect 1599 -45 1600 -44
rect 1604 -44 1612 -41
rect 1616 -38 1620 -37
rect 1604 -45 1605 -44
rect 1616 -49 1620 -42
rect 1583 -51 1620 -49
rect 1583 -53 1596 -51
rect 1600 -53 1620 -51
rect 1624 -48 1628 -30
rect 1624 -53 1628 -52
rect 1633 -28 1657 -16
rect 1637 -32 1657 -28
rect 1633 -37 1657 -32
rect 1633 -41 1653 -37
rect 1633 -53 1657 -41
rect 1662 -17 1666 -16
rect 1662 -39 1666 -21
rect 1670 -18 1690 -16
rect 1694 -18 1707 -16
rect 1670 -20 1707 -18
rect 1670 -27 1674 -20
rect 1685 -25 1686 -24
rect 1670 -32 1674 -31
rect 1678 -28 1686 -25
rect 1690 -25 1691 -24
rect 1690 -28 1699 -25
rect 1678 -29 1699 -28
rect 1678 -36 1682 -29
rect 1677 -37 1682 -36
rect 1662 -43 1671 -39
rect 1681 -41 1682 -37
rect 1677 -42 1682 -41
rect 1686 -34 1690 -33
rect 1667 -46 1671 -43
rect 1686 -46 1690 -38
rect 1667 -50 1690 -46
rect 1695 -45 1699 -29
rect 1703 -35 1707 -20
rect 1703 -40 1707 -39
rect 1713 -17 1721 10
rect 1731 -6 1747 -3
rect 1717 -21 1721 -17
rect 1713 -27 1727 -21
rect 1744 -25 1747 -6
rect 1785 -21 1791 171
rect 1713 -31 1723 -27
rect 1732 -26 1777 -25
rect 1732 -30 1735 -26
rect 1739 -29 1771 -26
rect 1739 -30 1740 -29
rect 1770 -30 1771 -29
rect 1775 -30 1777 -26
rect 1713 -35 1727 -31
rect 1713 -36 1739 -35
rect 1713 -40 1735 -36
rect 1713 -41 1739 -40
rect 1742 -37 1750 -33
rect 1754 -37 1769 -33
rect 1695 -49 1701 -45
rect 1705 -49 1706 -45
rect 1633 -57 1656 -53
rect 1660 -57 1663 -53
rect 1667 -57 1668 -53
rect 1582 -64 1609 -63
rect 1585 -67 1605 -64
rect 1614 -78 1628 -77
rect 1569 -83 1573 -79
rect 1589 -82 1590 -78
rect 1594 -82 1610 -78
rect 1614 -82 1615 -78
rect 1619 -82 1628 -78
rect 1569 -91 1577 -83
rect 1569 -92 1586 -91
rect 1569 -96 1582 -92
rect 1569 -97 1586 -96
rect 1590 -92 1596 -85
rect 1606 -86 1610 -82
rect 1622 -86 1623 -82
rect 1627 -86 1628 -82
rect 1606 -90 1609 -86
rect 1613 -90 1615 -86
rect 1622 -89 1628 -86
rect 1590 -94 1603 -92
rect 1452 -116 1523 -112
rect 1453 -146 1488 -142
rect 1435 -223 1459 -218
rect 1390 -236 1440 -232
rect 1390 -286 1394 -236
rect 1404 -240 1410 -236
rect 1414 -240 1440 -236
rect 1419 -245 1425 -240
rect 1419 -249 1420 -245
rect 1424 -249 1425 -245
rect 1431 -246 1436 -245
rect 1435 -250 1436 -246
rect 1431 -253 1436 -250
rect 1408 -257 1409 -253
rect 1413 -257 1428 -253
rect 1408 -262 1420 -261
rect 1408 -266 1412 -262
rect 1416 -266 1420 -262
rect 1408 -267 1420 -266
rect 1424 -262 1428 -257
rect 1435 -257 1436 -253
rect 1431 -258 1436 -257
rect 1405 -270 1412 -267
rect 1408 -275 1412 -270
rect 1424 -278 1428 -266
rect 1432 -278 1436 -258
rect 1408 -282 1409 -278
rect 1413 -282 1428 -278
rect 1431 -279 1436 -278
rect 1435 -283 1436 -279
rect 1431 -286 1436 -283
rect 1390 -289 1392 -286
rect 1423 -290 1431 -286
rect 1435 -290 1436 -286
rect 1423 -291 1436 -290
rect 1404 -300 1410 -296
rect 1414 -300 1420 -296
rect 1424 -300 1440 -296
rect 1404 -301 1440 -300
rect 1380 -304 1440 -301
rect 1305 -343 1308 -340
rect 1349 -343 1352 -326
rect 1359 -343 1362 -340
rect 1380 -343 1385 -304
rect 1432 -321 1435 -304
rect 1431 -325 1435 -321
rect 1406 -329 1442 -325
rect 1406 -333 1412 -329
rect 1416 -333 1422 -329
rect 1426 -333 1442 -329
rect 1425 -339 1438 -338
rect 1425 -343 1433 -339
rect 1437 -343 1438 -339
rect 1020 -346 1386 -343
rect 1036 -365 1039 -346
rect 1119 -348 1386 -346
rect 1433 -346 1438 -343
rect 1081 -363 1085 -361
rect 1119 -365 1122 -348
rect 1131 -355 1162 -352
rect 1081 -380 1085 -369
rect 1064 -384 1067 -381
rect 1081 -390 1084 -380
rect 1136 -385 1139 -382
rect 1081 -394 1082 -390
rect 1153 -391 1156 -369
rect 1159 -381 1162 -355
rect 1182 -365 1185 -348
rect 1192 -351 1195 -348
rect 1236 -365 1239 -348
rect 1246 -351 1249 -348
rect 1292 -365 1295 -348
rect 1302 -351 1305 -348
rect 1346 -365 1349 -348
rect 1356 -351 1359 -348
rect 1166 -374 1169 -369
rect 1199 -374 1202 -369
rect 1166 -377 1202 -374
rect 1159 -384 1164 -381
rect 1168 -385 1170 -382
rect 1190 -385 1191 -382
rect 1199 -386 1202 -377
rect 1220 -374 1223 -369
rect 1253 -374 1256 -369
rect 1220 -377 1256 -374
rect 1276 -374 1279 -369
rect 1309 -374 1312 -369
rect 1276 -377 1312 -374
rect 1206 -386 1209 -377
rect 1220 -382 1227 -381
rect 1220 -384 1224 -382
rect 1241 -386 1245 -383
rect 1199 -389 1209 -386
rect 1081 -402 1084 -394
rect 1153 -395 1154 -391
rect 1153 -403 1156 -395
rect 1199 -402 1202 -389
rect 1241 -390 1244 -386
rect 1253 -389 1256 -377
rect 1309 -378 1312 -377
rect 1319 -370 1321 -366
rect 1277 -385 1280 -382
rect 1253 -392 1272 -389
rect 1253 -402 1256 -392
rect 1301 -388 1304 -386
rect 1289 -396 1292 -390
rect 1303 -392 1304 -388
rect 1301 -393 1304 -392
rect 1266 -399 1292 -396
rect 1309 -402 1312 -382
rect 1047 -412 1050 -406
rect 1319 -405 1323 -370
rect 1330 -374 1333 -369
rect 1363 -374 1366 -369
rect 1330 -377 1366 -374
rect 1333 -386 1334 -383
rect 1352 -382 1358 -381
rect 1352 -384 1355 -382
rect 1333 -395 1336 -386
rect 1363 -387 1366 -377
rect 1335 -399 1336 -395
rect 1363 -402 1366 -391
rect 1119 -412 1122 -407
rect 1165 -412 1168 -406
rect 1219 -412 1222 -406
rect 1275 -412 1278 -406
rect 1322 -407 1323 -405
rect 1329 -412 1332 -406
rect 1012 -415 1366 -412
rect 1191 -418 1196 -415
rect 1297 -418 1301 -415
rect 667 -420 791 -419
rect 997 -422 1059 -418
rect 728 -431 1043 -426
rect 350 -446 356 -438
rect 350 -450 351 -446
rect 355 -450 356 -446
rect 361 -444 365 -443
rect 370 -444 376 -438
rect 411 -444 422 -441
rect 370 -448 371 -444
rect 375 -448 376 -444
rect 340 -451 345 -450
rect 340 -455 341 -451
rect 361 -451 365 -448
rect 340 -458 345 -455
rect 340 -462 341 -458
rect 340 -463 345 -462
rect 348 -455 361 -453
rect 348 -457 365 -455
rect 372 -455 403 -451
rect 340 -464 344 -463
rect 304 -468 344 -464
rect 301 -480 331 -477
rect 340 -481 344 -468
rect 348 -468 352 -457
rect 363 -464 368 -460
rect 372 -464 376 -455
rect 355 -472 358 -468
rect 362 -472 369 -468
rect 348 -476 352 -472
rect 348 -480 360 -476
rect 364 -477 369 -472
rect 340 -482 345 -481
rect 340 -486 341 -482
rect 345 -486 352 -483
rect 340 -489 352 -486
rect 356 -484 360 -480
rect 363 -481 379 -477
rect 356 -488 371 -484
rect 375 -488 376 -484
rect 399 -488 403 -455
rect 419 -454 422 -444
rect 443 -446 449 -438
rect 443 -450 444 -446
rect 448 -450 449 -446
rect 454 -444 458 -443
rect 463 -444 469 -438
rect 463 -448 464 -444
rect 468 -448 469 -444
rect 530 -446 536 -438
rect 509 -447 525 -446
rect 433 -451 438 -450
rect 433 -454 434 -451
rect 419 -455 434 -454
rect 454 -451 458 -448
rect 419 -457 438 -455
rect 433 -458 438 -457
rect 433 -462 434 -458
rect 433 -463 438 -462
rect 441 -455 454 -453
rect 441 -457 458 -455
rect 433 -481 437 -463
rect 441 -468 445 -457
rect 465 -460 469 -451
rect 513 -451 525 -447
rect 530 -450 531 -446
rect 535 -450 536 -446
rect 541 -444 545 -443
rect 550 -444 556 -438
rect 656 -441 1031 -438
rect 781 -442 1031 -441
rect 550 -448 551 -444
rect 555 -448 556 -444
rect 513 -452 521 -451
rect 520 -455 521 -452
rect 541 -451 545 -448
rect 520 -458 525 -455
rect 456 -464 461 -460
rect 465 -464 476 -460
rect 520 -462 521 -458
rect 520 -463 525 -462
rect 528 -455 541 -453
rect 528 -457 545 -455
rect 448 -472 451 -468
rect 455 -472 462 -468
rect 441 -476 445 -472
rect 441 -480 453 -476
rect 433 -482 438 -481
rect 433 -486 434 -482
rect 438 -486 445 -483
rect 433 -489 445 -486
rect 449 -484 453 -480
rect 457 -477 462 -472
rect 457 -481 472 -477
rect 520 -481 524 -463
rect 528 -468 532 -457
rect 552 -460 556 -451
rect 1002 -453 1005 -451
rect 1002 -456 1009 -453
rect 543 -464 548 -460
rect 552 -464 565 -460
rect 535 -472 538 -468
rect 542 -472 549 -468
rect 528 -476 532 -472
rect 528 -480 540 -476
rect 520 -482 525 -481
rect 449 -488 464 -484
rect 468 -488 469 -484
rect 520 -486 521 -482
rect 525 -486 532 -483
rect 520 -489 532 -486
rect 536 -484 540 -480
rect 544 -478 549 -472
rect 1002 -476 1005 -456
rect 544 -481 557 -478
rect 983 -477 1006 -476
rect 562 -481 1006 -477
rect 536 -488 551 -484
rect 555 -488 556 -484
rect 336 -498 342 -494
rect 346 -498 352 -494
rect 356 -498 380 -494
rect 429 -498 435 -494
rect 439 -498 445 -494
rect 449 -498 473 -494
rect 330 -499 473 -498
rect 516 -498 522 -494
rect 526 -498 532 -494
rect 536 -498 560 -494
rect 516 -499 560 -498
rect 330 -501 560 -499
rect 336 -502 380 -501
rect 429 -502 560 -501
rect 1025 -513 1030 -442
rect 1040 -500 1043 -431
rect 1055 -489 1059 -422
rect 1123 -421 1369 -418
rect 1123 -426 1126 -421
rect 1071 -431 1105 -427
rect 1169 -427 1172 -421
rect 1223 -427 1226 -421
rect 1279 -427 1282 -421
rect 1157 -438 1160 -430
rect 1157 -442 1158 -438
rect 1140 -451 1143 -448
rect 1157 -464 1160 -442
rect 1203 -444 1206 -431
rect 1203 -447 1213 -444
rect 1245 -447 1248 -443
rect 1257 -441 1260 -431
rect 1257 -444 1276 -441
rect 1305 -441 1308 -440
rect 1172 -451 1174 -448
rect 1194 -451 1195 -448
rect 1203 -456 1206 -447
rect 1170 -459 1206 -456
rect 1170 -464 1173 -459
rect 1203 -464 1206 -459
rect 1210 -456 1213 -447
rect 1224 -451 1228 -449
rect 1245 -450 1249 -447
rect 1224 -452 1231 -451
rect 1257 -456 1260 -444
rect 1307 -445 1308 -441
rect 1305 -447 1308 -445
rect 1281 -451 1284 -448
rect 1313 -451 1316 -431
rect 1313 -456 1316 -455
rect 1224 -459 1260 -456
rect 1224 -464 1227 -459
rect 1257 -464 1260 -459
rect 1280 -459 1316 -456
rect 1280 -464 1283 -459
rect 1313 -464 1316 -459
rect 1123 -487 1126 -468
rect 1186 -487 1189 -468
rect 1196 -487 1199 -482
rect 1240 -487 1243 -468
rect 1250 -487 1253 -482
rect 1296 -487 1299 -468
rect 1322 -479 1325 -428
rect 1333 -427 1336 -421
rect 1339 -438 1340 -434
rect 1337 -447 1340 -438
rect 1367 -442 1370 -431
rect 1337 -450 1338 -447
rect 1356 -451 1359 -449
rect 1356 -452 1362 -451
rect 1367 -456 1370 -446
rect 1334 -459 1370 -456
rect 1334 -464 1337 -459
rect 1367 -464 1370 -459
rect 1306 -487 1309 -482
rect 1350 -487 1353 -468
rect 1381 -479 1386 -348
rect 1410 -351 1411 -347
rect 1415 -351 1430 -347
rect 1437 -350 1438 -346
rect 1433 -351 1438 -350
rect 1404 -356 1415 -354
rect 1408 -360 1415 -356
rect 1410 -362 1415 -360
rect 1410 -363 1422 -362
rect 1410 -367 1414 -363
rect 1418 -367 1422 -363
rect 1410 -368 1422 -367
rect 1426 -363 1430 -351
rect 1426 -372 1430 -367
rect 1434 -371 1438 -351
rect 1410 -376 1411 -372
rect 1415 -376 1430 -372
rect 1433 -372 1438 -371
rect 1437 -376 1438 -372
rect 1433 -379 1438 -376
rect 1421 -384 1422 -380
rect 1426 -384 1427 -380
rect 1437 -383 1438 -379
rect 1433 -384 1438 -383
rect 1421 -389 1427 -384
rect 1406 -393 1412 -389
rect 1416 -393 1442 -389
rect 1406 -397 1442 -393
rect 1435 -411 1438 -397
rect 1408 -415 1444 -411
rect 1408 -419 1414 -415
rect 1418 -419 1444 -415
rect 1423 -424 1429 -419
rect 1423 -428 1424 -424
rect 1428 -428 1429 -424
rect 1435 -425 1440 -424
rect 1439 -429 1440 -425
rect 1435 -432 1440 -429
rect 1412 -436 1413 -432
rect 1417 -436 1432 -432
rect 1412 -441 1424 -440
rect 1412 -442 1416 -441
rect 1401 -445 1416 -442
rect 1420 -445 1424 -441
rect 1412 -446 1424 -445
rect 1428 -441 1432 -436
rect 1439 -436 1440 -432
rect 1435 -437 1440 -436
rect 1412 -454 1416 -446
rect 1428 -457 1432 -445
rect 1436 -457 1440 -437
rect 1412 -461 1413 -457
rect 1417 -461 1432 -457
rect 1435 -458 1440 -457
rect 1439 -462 1440 -458
rect 1435 -465 1440 -462
rect 1427 -469 1435 -465
rect 1439 -469 1440 -465
rect 1427 -470 1440 -469
rect 1454 -472 1459 -223
rect 1517 -230 1521 -116
rect 1547 -252 1550 -127
rect 1471 -256 1550 -252
rect 1569 -132 1577 -97
rect 1590 -98 1594 -94
rect 1598 -98 1603 -94
rect 1611 -103 1615 -90
rect 1633 -96 1657 -57
rect 1675 -63 1679 -50
rect 1713 -55 1727 -41
rect 1742 -46 1746 -37
rect 1757 -43 1761 -40
rect 1734 -50 1735 -46
rect 1739 -50 1746 -46
rect 1765 -41 1769 -37
rect 1773 -38 1777 -30
rect 1783 -27 1791 -21
rect 1787 -31 1791 -27
rect 1783 -37 1791 -31
rect 1780 -38 1791 -37
rect 1765 -45 1777 -41
rect 1784 -42 1791 -38
rect 1780 -43 1791 -42
rect 1749 -53 1753 -48
rect 1757 -49 1761 -47
rect 1757 -53 1770 -49
rect 1687 -59 1692 -55
rect 1696 -59 1700 -55
rect 1713 -56 1723 -55
rect 1687 -61 1700 -59
rect 1662 -71 1668 -64
rect 1675 -67 1677 -63
rect 1681 -67 1684 -63
rect 1680 -71 1684 -67
rect 1694 -68 1700 -61
rect 1704 -57 1723 -56
rect 1708 -59 1723 -57
rect 1727 -56 1739 -55
rect 1727 -59 1735 -56
rect 1708 -60 1735 -59
rect 1708 -61 1739 -60
rect 1748 -61 1758 -57
rect 1704 -62 1727 -61
rect 1713 -65 1727 -62
rect 1713 -70 1721 -65
rect 1767 -66 1770 -53
rect 1773 -56 1777 -45
rect 1773 -61 1777 -60
rect 1783 -65 1791 -43
rect 1662 -75 1671 -71
rect 1675 -75 1676 -71
rect 1680 -75 1696 -71
rect 1700 -75 1701 -71
rect 1717 -74 1721 -70
rect 1662 -76 1676 -75
rect 1672 -81 1675 -76
rect 1672 -84 1689 -81
rect 1622 -100 1623 -96
rect 1627 -100 1630 -96
rect 1634 -100 1657 -96
rect 1584 -108 1585 -104
rect 1589 -108 1595 -104
rect 1557 -249 1560 -134
rect 1569 -136 1573 -132
rect 1569 -149 1577 -136
rect 1583 -114 1587 -113
rect 1583 -133 1587 -118
rect 1591 -124 1595 -108
rect 1600 -107 1623 -103
rect 1600 -115 1604 -107
rect 1619 -110 1623 -107
rect 1600 -120 1604 -119
rect 1608 -112 1613 -111
rect 1608 -116 1609 -112
rect 1619 -114 1628 -110
rect 1608 -117 1613 -116
rect 1608 -124 1612 -117
rect 1591 -125 1612 -124
rect 1591 -128 1600 -125
rect 1599 -129 1600 -128
rect 1604 -128 1612 -125
rect 1616 -122 1620 -121
rect 1604 -129 1605 -128
rect 1616 -133 1620 -126
rect 1583 -137 1620 -133
rect 1624 -132 1628 -114
rect 1624 -137 1628 -136
rect 1633 -112 1657 -100
rect 1637 -116 1657 -112
rect 1633 -119 1657 -116
rect 1713 -91 1721 -74
rect 1633 -120 1674 -119
rect 1633 -124 1653 -120
rect 1657 -123 1674 -120
rect 1678 -123 1679 -119
rect 1686 -122 1689 -118
rect 1693 -122 1700 -118
rect 1695 -123 1700 -122
rect 1633 -134 1657 -124
rect 1606 -140 1610 -137
rect 1584 -144 1599 -141
rect 1633 -138 1653 -134
rect 1633 -142 1657 -138
rect 1662 -130 1663 -126
rect 1667 -130 1668 -126
rect 1699 -127 1700 -123
rect 1662 -132 1668 -130
rect 1662 -136 1663 -132
rect 1667 -133 1668 -132
rect 1678 -129 1691 -128
rect 1682 -133 1691 -129
rect 1695 -131 1700 -127
rect 1704 -120 1708 -119
rect 1667 -136 1675 -133
rect 1678 -134 1691 -133
rect 1704 -134 1708 -124
rect 1662 -139 1675 -136
rect 1687 -138 1708 -134
rect 1713 -138 1727 -91
rect 1745 -100 1780 -99
rect 1745 -104 1775 -100
rect 1678 -139 1682 -138
rect 1633 -143 1678 -142
rect 1596 -147 1599 -144
rect 1633 -146 1682 -143
rect 1687 -142 1691 -138
rect 1717 -142 1727 -138
rect 1569 -153 1573 -149
rect 1569 -159 1577 -153
rect 1582 -148 1620 -147
rect 1582 -152 1585 -148
rect 1589 -151 1608 -148
rect 1589 -152 1590 -151
rect 1607 -152 1608 -151
rect 1612 -151 1620 -148
rect 1633 -148 1657 -146
rect 1687 -147 1691 -146
rect 1633 -149 1653 -148
rect 1612 -152 1613 -151
rect 1582 -159 1588 -152
rect 1637 -152 1653 -149
rect 1702 -149 1708 -142
rect 1677 -150 1678 -149
rect 1637 -153 1657 -152
rect 1599 -155 1603 -154
rect 1633 -155 1657 -153
rect 1670 -153 1678 -150
rect 1682 -150 1683 -149
rect 1700 -150 1701 -149
rect 1682 -153 1691 -150
rect 1670 -154 1691 -153
rect 1695 -153 1701 -150
rect 1705 -153 1708 -149
rect 1695 -154 1708 -153
rect 1713 -147 1727 -142
rect 1713 -148 1767 -147
rect 1717 -152 1767 -148
rect 1713 -155 1727 -152
rect 1569 -163 1573 -159
rect 1599 -163 1603 -159
rect 1608 -158 1657 -155
rect 1612 -159 1657 -158
rect 1608 -163 1612 -162
rect 1569 -187 1577 -163
rect 1582 -167 1603 -163
rect 1615 -165 1628 -162
rect 1582 -177 1586 -167
rect 1599 -168 1612 -167
rect 1615 -168 1623 -165
rect 1582 -182 1586 -181
rect 1590 -174 1595 -170
rect 1599 -172 1608 -168
rect 1599 -173 1612 -172
rect 1622 -169 1623 -168
rect 1627 -169 1628 -165
rect 1622 -171 1628 -169
rect 1590 -178 1591 -174
rect 1622 -175 1623 -171
rect 1627 -175 1628 -171
rect 1633 -163 1657 -159
rect 1637 -167 1657 -163
rect 1633 -177 1657 -167
rect 1717 -169 1727 -155
rect 1717 -172 1719 -169
rect 1590 -179 1595 -178
rect 1590 -183 1598 -179
rect 1602 -183 1604 -179
rect 1611 -182 1612 -178
rect 1616 -181 1633 -178
rect 1637 -180 1657 -177
rect 1637 -181 1641 -180
rect 1616 -182 1641 -181
rect 1633 -186 1641 -182
rect 1647 -184 1657 -180
rect 1788 -184 1792 -65
rect 1647 -186 1792 -184
rect 1633 -187 1792 -186
rect 1571 -215 1576 -187
rect 1649 -188 1792 -187
rect 1768 -189 1792 -188
rect 1672 -200 1715 -195
rect 1766 -197 1771 -196
rect 1571 -216 1697 -215
rect 1571 -221 1692 -216
rect 1641 -234 1642 -232
rect 1728 -230 1729 -227
rect 1733 -230 1758 -227
rect 1641 -238 1647 -234
rect 1641 -243 1649 -238
rect 1705 -239 1713 -238
rect 1766 -239 1771 -202
rect 1641 -244 1666 -243
rect 1641 -248 1645 -244
rect 1649 -247 1666 -244
rect 1670 -247 1671 -243
rect 1678 -246 1680 -242
rect 1684 -246 1692 -242
rect 1687 -247 1692 -246
rect 1557 -259 1561 -249
rect 1641 -258 1649 -248
rect 1641 -262 1645 -258
rect 1641 -266 1649 -262
rect 1654 -254 1655 -250
rect 1659 -254 1660 -250
rect 1691 -251 1692 -247
rect 1654 -256 1660 -254
rect 1654 -260 1655 -256
rect 1659 -257 1660 -256
rect 1670 -253 1683 -252
rect 1674 -257 1683 -253
rect 1687 -255 1692 -251
rect 1696 -244 1700 -243
rect 1659 -260 1667 -257
rect 1670 -258 1683 -257
rect 1696 -258 1700 -248
rect 1654 -263 1667 -260
rect 1679 -262 1700 -258
rect 1705 -244 1771 -239
rect 1705 -262 1713 -244
rect 1670 -263 1674 -262
rect 1641 -267 1670 -266
rect 1641 -270 1674 -267
rect 1679 -266 1683 -262
rect 1709 -266 1713 -262
rect 1641 -272 1649 -270
rect 1679 -271 1683 -270
rect 1641 -276 1645 -272
rect 1694 -273 1700 -266
rect 1669 -274 1670 -273
rect 1641 -309 1649 -276
rect 1662 -277 1670 -274
rect 1674 -274 1675 -273
rect 1692 -274 1693 -273
rect 1674 -277 1693 -274
rect 1697 -277 1700 -273
rect 1662 -278 1700 -277
rect 1705 -272 1713 -266
rect 1709 -276 1713 -272
rect 1683 -281 1686 -278
rect 1683 -284 1698 -281
rect 1668 -288 1671 -285
rect 1641 -313 1645 -309
rect 1641 -325 1649 -313
rect 1654 -289 1658 -288
rect 1654 -311 1658 -293
rect 1662 -292 1699 -288
rect 1662 -299 1666 -292
rect 1677 -297 1678 -296
rect 1662 -304 1666 -303
rect 1670 -300 1678 -297
rect 1682 -297 1683 -296
rect 1682 -300 1691 -297
rect 1670 -301 1691 -300
rect 1670 -308 1674 -301
rect 1669 -309 1674 -308
rect 1654 -315 1663 -311
rect 1673 -313 1674 -309
rect 1669 -314 1674 -313
rect 1678 -306 1682 -305
rect 1659 -318 1663 -315
rect 1678 -318 1682 -310
rect 1659 -322 1682 -318
rect 1687 -317 1691 -301
rect 1695 -307 1699 -292
rect 1695 -312 1699 -311
rect 1705 -289 1713 -276
rect 1709 -293 1713 -289
rect 1687 -321 1693 -317
rect 1697 -321 1698 -317
rect 1641 -329 1648 -325
rect 1652 -329 1655 -325
rect 1659 -329 1660 -325
rect 1641 -393 1649 -329
rect 1667 -335 1671 -322
rect 1679 -331 1684 -327
rect 1688 -331 1692 -327
rect 1705 -328 1713 -293
rect 1730 -308 1734 -267
rect 1815 -273 1818 503
rect 1829 199 1834 502
rect 1829 198 1835 199
rect 1779 -276 1819 -273
rect 1741 -293 1794 -292
rect 1830 -293 1835 198
rect 1741 -295 1835 -293
rect 1778 -297 1835 -295
rect 1830 -298 1835 -297
rect 1730 -313 1741 -308
rect 1679 -333 1692 -331
rect 1654 -339 1660 -336
rect 1667 -339 1669 -335
rect 1673 -339 1676 -335
rect 1654 -343 1655 -339
rect 1659 -343 1660 -339
rect 1672 -343 1676 -339
rect 1686 -340 1692 -333
rect 1696 -329 1713 -328
rect 1700 -333 1713 -329
rect 1696 -334 1713 -333
rect 1705 -342 1713 -334
rect 1654 -347 1663 -343
rect 1667 -347 1668 -343
rect 1672 -347 1688 -343
rect 1692 -347 1693 -343
rect 1709 -346 1713 -342
rect 1654 -348 1668 -347
rect 1655 -360 1658 -348
rect 1655 -363 1698 -360
rect 1641 -397 1645 -393
rect 1641 -409 1649 -397
rect 1654 -373 1658 -372
rect 1654 -395 1658 -377
rect 1662 -374 1682 -372
rect 1686 -374 1699 -372
rect 1662 -376 1699 -374
rect 1662 -383 1666 -376
rect 1677 -381 1678 -380
rect 1662 -388 1666 -387
rect 1670 -384 1678 -381
rect 1682 -381 1683 -380
rect 1682 -384 1691 -381
rect 1670 -385 1691 -384
rect 1670 -392 1674 -385
rect 1669 -393 1674 -392
rect 1654 -399 1663 -395
rect 1673 -397 1674 -393
rect 1669 -398 1674 -397
rect 1678 -390 1682 -389
rect 1659 -402 1663 -399
rect 1678 -402 1682 -394
rect 1659 -406 1682 -402
rect 1687 -401 1691 -385
rect 1695 -391 1699 -376
rect 1695 -396 1699 -395
rect 1705 -373 1713 -346
rect 1719 -338 1725 -335
rect 1719 -370 1722 -338
rect 1709 -377 1713 -373
rect 1705 -383 1719 -377
rect 1736 -381 1741 -313
rect 1705 -387 1715 -383
rect 1724 -382 1769 -381
rect 1724 -386 1727 -382
rect 1731 -385 1763 -382
rect 1731 -386 1732 -385
rect 1762 -386 1763 -385
rect 1767 -386 1769 -382
rect 1705 -391 1719 -387
rect 1705 -392 1731 -391
rect 1705 -396 1727 -392
rect 1705 -397 1731 -396
rect 1734 -393 1742 -389
rect 1746 -393 1761 -389
rect 1687 -405 1693 -401
rect 1697 -405 1698 -401
rect 1641 -413 1648 -409
rect 1652 -413 1655 -409
rect 1659 -413 1660 -409
rect 1408 -479 1414 -475
rect 1418 -479 1424 -475
rect 1428 -479 1444 -475
rect 1641 -475 1649 -413
rect 1667 -419 1671 -406
rect 1705 -411 1719 -397
rect 1734 -402 1738 -393
rect 1749 -399 1753 -396
rect 1726 -406 1727 -402
rect 1731 -406 1738 -402
rect 1757 -397 1761 -393
rect 1765 -394 1769 -386
rect 1775 -383 1783 -377
rect 1779 -387 1783 -383
rect 1775 -393 1783 -387
rect 1772 -394 1783 -393
rect 1757 -401 1769 -397
rect 1776 -398 1783 -394
rect 1772 -399 1783 -398
rect 1741 -409 1745 -404
rect 1749 -405 1753 -403
rect 1749 -409 1762 -405
rect 1679 -415 1684 -411
rect 1688 -415 1692 -411
rect 1705 -412 1715 -411
rect 1679 -417 1692 -415
rect 1654 -427 1660 -420
rect 1667 -423 1669 -419
rect 1673 -423 1676 -419
rect 1686 -421 1692 -417
rect 1696 -413 1715 -412
rect 1700 -415 1715 -413
rect 1719 -412 1731 -411
rect 1719 -415 1727 -412
rect 1700 -416 1727 -415
rect 1700 -417 1731 -416
rect 1734 -413 1737 -410
rect 1759 -413 1762 -409
rect 1738 -417 1750 -413
rect 1758 -417 1762 -413
rect 1765 -412 1769 -401
rect 1765 -417 1769 -416
rect 1696 -418 1719 -417
rect 1672 -427 1676 -423
rect 1686 -424 1701 -421
rect 1654 -431 1663 -427
rect 1667 -431 1668 -427
rect 1672 -431 1688 -427
rect 1692 -431 1693 -427
rect 1654 -432 1668 -431
rect 1664 -437 1667 -432
rect 1664 -440 1681 -437
rect 1698 -448 1701 -424
rect 1705 -425 1713 -418
rect 1775 -421 1783 -399
rect 1831 -411 1835 -310
rect 1831 -414 1836 -411
rect 1725 -425 1734 -422
rect 1747 -425 1769 -422
rect 1780 -425 1784 -421
rect 1705 -426 1718 -425
rect 1709 -430 1718 -426
rect 1731 -429 1734 -425
rect 1705 -440 1718 -430
rect 1723 -430 1763 -429
rect 1723 -434 1724 -430
rect 1728 -433 1752 -430
rect 1728 -434 1729 -433
rect 1751 -434 1752 -433
rect 1756 -434 1759 -430
rect 1733 -437 1737 -436
rect 1705 -444 1720 -440
rect 1724 -444 1725 -440
rect 1766 -439 1769 -425
rect 1641 -476 1666 -475
rect 1360 -487 1363 -482
rect 1381 -483 1444 -479
rect 1641 -480 1645 -476
rect 1649 -479 1666 -476
rect 1670 -479 1671 -475
rect 1678 -478 1681 -474
rect 1685 -478 1692 -474
rect 1687 -479 1692 -478
rect 1381 -487 1386 -483
rect 1121 -490 1386 -487
rect 1641 -490 1649 -480
rect 1641 -494 1645 -490
rect 1641 -498 1649 -494
rect 1654 -486 1655 -482
rect 1659 -486 1660 -482
rect 1691 -483 1692 -479
rect 1654 -488 1660 -486
rect 1654 -492 1655 -488
rect 1659 -489 1660 -488
rect 1670 -485 1683 -484
rect 1674 -489 1683 -485
rect 1687 -487 1692 -483
rect 1696 -476 1700 -475
rect 1659 -492 1667 -489
rect 1670 -490 1683 -489
rect 1696 -490 1700 -480
rect 1654 -495 1667 -492
rect 1679 -494 1700 -490
rect 1705 -494 1718 -444
rect 1723 -450 1727 -449
rect 1733 -450 1737 -441
rect 1774 -440 1784 -425
rect 1772 -441 1784 -440
rect 1742 -447 1743 -443
rect 1747 -446 1760 -443
rect 1776 -445 1784 -441
rect 1772 -446 1784 -445
rect 1747 -447 1764 -446
rect 1756 -449 1764 -447
rect 1723 -470 1727 -454
rect 1731 -454 1752 -450
rect 1731 -460 1735 -454
rect 1748 -457 1752 -454
rect 1756 -457 1757 -453
rect 1731 -465 1735 -464
rect 1739 -461 1740 -457
rect 1744 -460 1745 -457
rect 1744 -461 1752 -460
rect 1739 -465 1752 -461
rect 1760 -465 1764 -449
rect 1723 -474 1724 -470
rect 1728 -474 1731 -470
rect 1735 -474 1736 -470
rect 1740 -476 1744 -472
rect 1724 -480 1728 -479
rect 1731 -480 1740 -477
rect 1731 -481 1744 -480
rect 1724 -485 1728 -484
rect 1740 -483 1744 -481
rect 1724 -489 1736 -485
rect 1670 -495 1674 -494
rect 1040 -501 1435 -500
rect 1040 -505 1583 -501
rect 1641 -499 1670 -498
rect 1641 -502 1674 -499
rect 1679 -498 1683 -494
rect 1709 -496 1718 -494
rect 1709 -497 1721 -496
rect 1709 -498 1717 -497
rect 1612 -507 1631 -504
rect 1641 -504 1649 -502
rect 1679 -503 1683 -502
rect 1641 -508 1645 -504
rect 1694 -505 1700 -498
rect 1669 -506 1670 -505
rect 1295 -513 1630 -512
rect 1025 -515 1631 -513
rect 1025 -516 1308 -515
rect 1313 -524 1352 -523
rect 1518 -524 1607 -522
rect 1313 -528 1607 -524
rect 1612 -528 1613 -522
rect 949 -540 1485 -536
rect 1153 -541 1485 -540
rect 1113 -550 1581 -549
rect 1020 -553 1581 -550
rect 1020 -554 1299 -553
rect 1575 -554 1581 -553
rect 1020 -555 1127 -554
rect 1575 -555 1578 -554
rect 1360 -566 1473 -562
rect 1360 -567 1480 -566
rect 1627 -581 1631 -515
rect 1641 -540 1649 -508
rect 1662 -509 1670 -506
rect 1674 -506 1675 -505
rect 1692 -506 1693 -505
rect 1674 -509 1683 -506
rect 1662 -510 1683 -509
rect 1687 -509 1693 -506
rect 1697 -509 1700 -505
rect 1687 -510 1700 -509
rect 1705 -501 1717 -498
rect 1705 -502 1721 -501
rect 1724 -497 1728 -492
rect 1705 -504 1718 -502
rect 1709 -508 1718 -504
rect 1705 -511 1718 -508
rect 1710 -525 1718 -511
rect 1724 -508 1728 -501
rect 1732 -501 1736 -489
rect 1740 -490 1744 -487
rect 1748 -493 1752 -465
rect 1739 -497 1740 -493
rect 1744 -497 1752 -493
rect 1748 -498 1752 -497
rect 1756 -469 1764 -465
rect 1756 -488 1760 -469
rect 1774 -475 1784 -446
rect 1764 -476 1784 -475
rect 1768 -480 1771 -476
rect 1775 -480 1784 -476
rect 1764 -481 1784 -480
rect 1760 -492 1763 -488
rect 1767 -492 1768 -488
rect 1756 -501 1760 -492
rect 1774 -497 1784 -481
rect 1732 -503 1760 -501
rect 1764 -498 1784 -497
rect 1768 -502 1771 -498
rect 1775 -502 1784 -498
rect 1764 -503 1784 -502
rect 1732 -505 1740 -503
rect 1739 -507 1740 -505
rect 1744 -505 1760 -503
rect 1744 -507 1745 -505
rect 1748 -510 1749 -508
rect 1728 -512 1749 -510
rect 1753 -512 1756 -508
rect 1760 -512 1761 -508
rect 1724 -514 1761 -512
rect 1774 -525 1784 -503
rect 1658 -532 1692 -528
rect 1780 -540 1784 -525
rect 1641 -544 1784 -540
rect 1760 -545 1784 -544
rect 1659 -554 1674 -550
rect 1697 -550 1749 -547
rect 1832 -549 1836 -414
rect 1756 -550 1836 -549
rect 1645 -566 1704 -562
rect 1663 -581 1667 -576
rect 1699 -575 1704 -566
rect 1731 -569 1734 -558
rect 1745 -562 1749 -550
rect 1759 -553 1836 -550
rect 1745 -565 1794 -562
rect 1718 -572 1769 -569
rect 1699 -581 1806 -575
rect 1627 -584 1667 -581
<< metal2 >>
rect 1457 537 1463 538
rect 1456 536 1559 537
rect 1840 536 1844 537
rect 1456 532 1844 536
rect 499 480 850 481
rect 1457 480 1463 532
rect 1555 531 1844 532
rect 1772 497 1775 503
rect 499 476 1463 480
rect 363 455 468 456
rect 363 453 463 455
rect 81 448 110 452
rect 17 444 84 448
rect 17 302 22 444
rect 91 437 344 441
rect 32 379 36 430
rect 91 402 96 437
rect 339 433 343 437
rect 109 424 110 427
rect 114 424 198 427
rect 202 424 291 427
rect 295 424 316 427
rect 313 421 316 424
rect 363 421 367 453
rect 467 453 468 455
rect 413 441 416 442
rect 413 438 462 441
rect 413 422 416 438
rect 474 423 478 457
rect 499 441 504 476
rect 846 475 1463 476
rect 1457 474 1463 475
rect 945 450 946 455
rect 503 437 504 441
rect 516 438 764 442
rect 516 434 520 438
rect 573 426 662 429
rect 571 425 662 426
rect 666 425 749 429
rect 313 417 367 421
rect 195 406 339 409
rect 521 408 668 411
rect 90 398 102 402
rect 195 402 198 406
rect 665 404 668 408
rect 107 398 118 402
rect 247 397 248 400
rect 31 377 36 379
rect 31 341 35 377
rect 175 376 223 379
rect 175 375 232 376
rect 220 372 232 375
rect 245 366 248 397
rect 288 392 291 398
rect 569 400 573 403
rect 288 389 339 392
rect 569 392 572 400
rect 521 389 572 392
rect 665 400 666 404
rect 683 402 702 406
rect 760 404 764 438
rect 945 414 949 450
rect 1003 441 1025 444
rect 981 414 984 437
rect 1090 424 1170 427
rect 1090 418 1093 424
rect 1051 415 1093 418
rect 1166 418 1169 424
rect 1190 422 1249 425
rect 981 411 996 414
rect 1123 414 1144 417
rect 746 400 754 404
rect 759 402 764 404
rect 759 400 986 402
rect 566 381 569 389
rect 493 378 504 380
rect 566 378 580 381
rect 493 377 498 378
rect 274 374 498 377
rect 502 374 504 378
rect 274 373 504 374
rect 604 372 607 399
rect 666 390 669 400
rect 760 399 986 400
rect 773 398 986 399
rect 972 390 976 391
rect 666 386 976 390
rect 619 378 678 381
rect 509 369 607 372
rect 706 378 968 381
rect 692 374 696 377
rect 692 371 759 374
rect 197 365 250 366
rect 115 362 250 365
rect 509 364 513 369
rect 115 356 118 362
rect 64 353 129 356
rect 31 337 72 341
rect 68 330 72 337
rect 21 298 22 302
rect 29 328 32 329
rect 29 325 36 328
rect 29 260 32 325
rect 72 326 105 329
rect 125 329 128 353
rect 207 353 292 356
rect 296 353 318 356
rect 393 355 458 358
rect 265 343 307 346
rect 315 336 318 353
rect 454 352 458 355
rect 509 352 512 364
rect 755 361 759 371
rect 516 358 536 360
rect 516 357 532 358
rect 516 353 517 357
rect 521 354 532 357
rect 536 355 621 358
rect 720 358 785 361
rect 521 353 536 354
rect 516 352 524 353
rect 351 346 418 349
rect 326 343 354 346
rect 454 349 512 352
rect 314 332 318 336
rect 176 325 209 328
rect 189 321 192 325
rect 301 321 304 327
rect 189 318 304 321
rect 265 309 266 312
rect 263 261 266 309
rect 314 303 317 332
rect 358 327 365 330
rect 308 299 342 303
rect 302 298 342 299
rect 29 257 123 260
rect 133 258 276 261
rect 120 253 123 257
rect 271 227 302 231
rect 252 226 276 227
rect 209 223 276 226
rect 209 222 212 223
rect 153 219 212 222
rect 153 210 157 219
rect 315 212 318 298
rect 326 275 347 279
rect 358 262 361 327
rect 401 328 434 331
rect 454 331 457 349
rect 593 347 751 350
rect 409 314 410 319
rect 409 271 412 314
rect 419 279 423 328
rect 505 327 538 330
rect 518 323 521 327
rect 630 323 633 329
rect 518 320 633 323
rect 685 330 692 333
rect 594 311 595 314
rect 509 290 512 291
rect 509 287 579 290
rect 509 278 512 287
rect 457 275 512 278
rect 457 271 460 275
rect 409 268 461 271
rect 592 263 595 311
rect 635 301 669 305
rect 629 300 669 301
rect 645 272 673 275
rect 685 265 688 330
rect 728 331 761 334
rect 781 334 784 358
rect 863 358 948 361
rect 840 350 914 352
rect 840 349 918 350
rect 744 276 748 331
rect 832 330 865 333
rect 845 326 848 330
rect 957 326 960 332
rect 845 323 960 326
rect 753 289 756 314
rect 921 314 922 317
rect 770 277 829 280
rect 837 276 841 314
rect 919 266 922 314
rect 358 259 452 262
rect 462 260 605 263
rect 685 262 779 265
rect 789 263 932 266
rect 449 255 452 259
rect 776 258 779 262
rect 747 251 767 254
rect 747 249 750 251
rect 507 246 750 249
rect 764 250 767 251
rect 827 251 875 254
rect 764 246 766 250
rect 770 246 771 249
rect 507 230 510 246
rect 827 242 830 251
rect 758 240 830 242
rect 754 239 830 240
rect 836 233 841 236
rect 327 227 510 230
rect 536 229 841 233
rect 536 228 659 229
rect 537 212 542 228
rect 869 215 872 251
rect 63 207 157 210
rect 28 179 35 182
rect 28 114 31 179
rect 71 180 104 183
rect 124 183 127 207
rect 206 207 291 210
rect 315 209 319 212
rect 261 198 308 201
rect 261 191 264 198
rect 316 192 319 209
rect 392 209 457 212
rect 315 189 319 192
rect 424 193 427 209
rect 85 145 88 180
rect 175 179 208 182
rect 188 175 191 179
rect 300 175 303 181
rect 188 172 303 175
rect 264 163 265 166
rect 185 147 188 163
rect 85 141 178 145
rect 184 144 251 147
rect 173 128 178 141
rect 173 124 246 128
rect 262 115 265 163
rect 315 159 318 189
rect 357 181 364 184
rect 310 158 340 159
rect 310 153 339 158
rect 280 124 300 128
rect 28 111 122 114
rect 132 112 275 115
rect 119 107 122 111
rect 181 0 182 4
rect 311 10 317 153
rect 325 144 348 147
rect 338 128 342 129
rect 326 124 342 128
rect 338 103 342 124
rect 357 116 360 181
rect 400 182 433 185
rect 453 185 456 209
rect 535 209 620 212
rect 719 212 784 215
rect 668 204 679 205
rect 590 201 679 204
rect 590 197 593 201
rect 415 135 418 182
rect 504 181 537 184
rect 517 177 520 181
rect 629 177 632 183
rect 517 174 632 177
rect 675 171 678 201
rect 684 184 691 187
rect 424 169 427 170
rect 593 165 594 168
rect 674 167 680 171
rect 424 143 427 165
rect 415 131 514 135
rect 591 117 594 165
rect 633 155 669 158
rect 607 131 666 136
rect 357 113 451 116
rect 461 114 604 117
rect 448 109 451 113
rect 338 99 415 103
rect 412 95 415 99
rect 495 98 497 103
rect 495 95 500 98
rect 370 91 383 94
rect 370 81 373 91
rect 370 78 385 81
rect 396 66 400 91
rect 412 91 500 95
rect 412 90 415 91
rect 411 77 585 80
rect 677 75 680 167
rect 684 119 687 184
rect 727 185 760 188
rect 780 188 783 212
rect 862 212 947 215
rect 955 206 958 236
rect 925 203 958 206
rect 925 198 929 203
rect 920 195 929 198
rect 747 149 751 185
rect 831 184 864 187
rect 844 180 847 184
rect 956 180 959 186
rect 844 177 959 180
rect 920 168 921 171
rect 731 145 751 149
rect 747 144 751 145
rect 705 133 832 136
rect 838 133 839 136
rect 705 132 839 133
rect 918 120 921 168
rect 684 116 778 119
rect 788 117 931 120
rect 775 112 778 116
rect 727 108 731 109
rect 727 59 731 104
rect 965 98 968 378
rect 502 56 731 59
rect 502 55 727 56
rect 964 46 968 98
rect 469 42 503 46
rect 558 43 968 46
rect 964 42 968 43
rect 499 38 503 42
rect 499 35 568 38
rect 565 31 568 35
rect 972 31 976 386
rect 373 25 461 29
rect 466 25 546 28
rect 565 27 976 31
rect 983 17 986 398
rect 993 302 996 411
rect 1127 408 1130 414
rect 1170 414 1196 417
rect 1200 414 1201 417
rect 1246 416 1249 422
rect 1270 417 1289 420
rect 1246 413 1253 416
rect 1270 412 1273 417
rect 1293 418 1332 419
rect 1293 416 1328 418
rect 1120 407 1130 408
rect 1156 407 1175 410
rect 1066 404 1078 407
rect 1120 405 1122 407
rect 1075 340 1078 404
rect 1126 405 1130 407
rect 1138 404 1159 407
rect 1172 404 1220 407
rect 1283 407 1342 410
rect 1253 402 1256 405
rect 1163 387 1166 399
rect 1088 384 1166 387
rect 1253 399 1311 402
rect 1088 355 1091 384
rect 1242 380 1246 398
rect 1123 376 1246 380
rect 1123 350 1127 376
rect 1242 375 1246 376
rect 1257 361 1315 364
rect 1142 356 1224 359
rect 1257 358 1260 361
rect 1287 353 1346 356
rect 1127 346 1148 349
rect 1174 346 1200 349
rect 1204 346 1205 349
rect 1250 347 1257 350
rect 1170 340 1173 346
rect 1075 337 1173 340
rect 1250 341 1253 347
rect 1297 345 1332 347
rect 1297 344 1336 345
rect 1194 338 1253 341
rect 1089 317 1161 319
rect 1085 315 1161 317
rect 993 299 1108 302
rect 993 298 1006 299
rect 1157 282 1161 315
rect 1303 308 1306 344
rect 1433 308 1443 309
rect 1303 305 1374 308
rect 1090 279 1170 282
rect 1370 281 1373 305
rect 1433 307 1435 308
rect 1426 303 1435 307
rect 1440 303 1443 308
rect 1426 302 1443 303
rect 1090 273 1093 279
rect 1051 270 1093 273
rect 1166 272 1169 279
rect 1190 277 1249 280
rect 1051 228 1054 270
rect 1123 269 1144 272
rect 1170 269 1196 272
rect 1200 269 1201 272
rect 1246 271 1249 277
rect 1270 272 1289 275
rect 1246 268 1253 271
rect 1270 267 1273 272
rect 1293 273 1332 274
rect 1293 271 1328 273
rect 1066 259 1078 262
rect 1050 162 1054 228
rect 1075 195 1078 259
rect 1138 259 1220 262
rect 1283 262 1342 265
rect 1253 257 1256 260
rect 1253 254 1311 257
rect 1242 235 1246 253
rect 1352 239 1369 242
rect 1431 236 1477 239
rect 1123 231 1246 235
rect 1123 205 1127 231
rect 1242 230 1246 231
rect 1257 216 1315 219
rect 1142 211 1224 214
rect 1257 213 1260 216
rect 1287 208 1346 211
rect 1474 206 1477 236
rect 1489 221 1493 485
rect 1507 343 1510 495
rect 1644 494 1775 497
rect 1559 467 1562 494
rect 1526 449 1597 452
rect 1526 361 1529 449
rect 1594 445 1597 449
rect 1522 358 1529 361
rect 1541 396 1580 400
rect 1507 340 1515 343
rect 1512 335 1515 340
rect 1512 332 1522 335
rect 1519 311 1522 332
rect 1514 285 1520 290
rect 1514 280 1515 285
rect 1514 279 1520 280
rect 1489 218 1523 221
rect 1481 206 1510 207
rect 1127 201 1148 204
rect 1174 201 1200 204
rect 1204 201 1205 204
rect 1250 202 1257 205
rect 1170 195 1173 201
rect 1075 192 1173 195
rect 1250 196 1253 202
rect 1297 200 1332 202
rect 1474 203 1510 206
rect 1336 200 1372 202
rect 1297 199 1372 200
rect 1425 202 1429 203
rect 1408 199 1433 202
rect 1194 193 1253 196
rect 1340 171 1344 174
rect 999 154 1046 157
rect 392 14 986 17
rect 289 5 312 10
rect 285 3 312 5
rect 181 -20 185 0
rect 181 -21 552 -20
rect 181 -22 921 -21
rect 181 -24 976 -22
rect 181 -25 185 -24
rect 550 -25 976 -24
rect 908 -26 976 -25
rect 20 -39 370 -36
rect 92 -58 121 -54
rect 28 -62 95 -58
rect 28 -105 33 -62
rect 102 -69 355 -65
rect -8 -110 33 -105
rect 28 -204 33 -110
rect 43 -127 47 -76
rect 102 -104 107 -69
rect 350 -73 354 -69
rect 120 -82 121 -79
rect 125 -82 209 -79
rect 213 -82 302 -79
rect 206 -100 350 -97
rect 101 -108 113 -104
rect 206 -104 209 -100
rect 118 -108 129 -104
rect 258 -109 259 -106
rect 42 -129 47 -127
rect 42 -165 46 -129
rect 186 -130 234 -127
rect 186 -131 243 -130
rect 231 -134 243 -131
rect 256 -140 259 -109
rect 299 -114 302 -108
rect 299 -117 350 -114
rect 365 -117 370 -39
rect 392 -104 395 -35
rect 411 -93 414 -35
rect 423 -71 426 -35
rect 435 -87 436 -82
rect 485 -83 489 -49
rect 527 -68 775 -64
rect 527 -72 531 -68
rect 535 -80 580 -79
rect 584 -80 673 -77
rect 499 -81 502 -80
rect 432 -106 436 -87
rect 497 -84 502 -81
rect 535 -81 673 -80
rect 677 -81 760 -77
rect 535 -82 583 -81
rect 535 -84 538 -82
rect 497 -87 538 -84
rect 432 -109 486 -106
rect 497 -117 502 -87
rect 532 -98 679 -95
rect 676 -102 679 -98
rect 524 -104 531 -103
rect 524 -106 525 -104
rect 518 -108 525 -106
rect 529 -108 531 -104
rect 518 -109 531 -108
rect 580 -106 584 -103
rect 580 -114 583 -106
rect 532 -117 583 -114
rect 676 -106 677 -102
rect 694 -104 713 -100
rect 771 -102 775 -68
rect 991 -90 994 34
rect 999 30 1002 154
rect 1043 153 1046 154
rect 1062 154 1105 157
rect 1109 154 1110 157
rect 1062 153 1065 154
rect 1043 150 1065 153
rect 1089 137 1169 140
rect 1089 131 1092 137
rect 1050 128 1092 131
rect 1165 130 1168 137
rect 1189 135 1248 138
rect 1417 136 1420 137
rect 1122 127 1143 130
rect 1169 127 1195 130
rect 1199 127 1200 130
rect 1245 129 1248 135
rect 1269 130 1288 133
rect 1245 126 1252 129
rect 1269 125 1272 130
rect 1407 133 1420 136
rect 1292 131 1331 132
rect 1292 129 1327 131
rect 1353 127 1372 130
rect 1065 117 1077 120
rect 1074 53 1077 117
rect 1137 117 1219 120
rect 1282 120 1341 123
rect 1252 115 1255 118
rect 1252 112 1310 115
rect 1241 93 1245 111
rect 1122 89 1245 93
rect 1122 63 1126 89
rect 1241 88 1245 89
rect 1256 74 1314 77
rect 1141 69 1223 72
rect 1256 71 1259 74
rect 1286 66 1345 69
rect 1126 59 1147 62
rect 1173 59 1199 62
rect 1203 59 1204 62
rect 1249 60 1256 63
rect 1169 53 1172 59
rect 1011 49 1063 51
rect 1074 50 1172 53
rect 1249 54 1252 60
rect 1296 58 1331 60
rect 1353 60 1356 127
rect 1335 58 1356 60
rect 1296 57 1356 58
rect 1360 91 1395 95
rect 1193 51 1252 54
rect 1011 48 1059 49
rect 1299 43 1306 44
rect 1299 41 1300 43
rect 1015 38 1300 41
rect 1305 38 1306 43
rect 1299 37 1306 38
rect 1013 33 1020 34
rect 1013 28 1014 33
rect 1019 30 1058 33
rect 1360 33 1363 91
rect 1417 87 1420 133
rect 1369 83 1420 87
rect 1019 28 1020 30
rect 1096 29 1353 32
rect 1357 30 1365 33
rect 1013 27 1020 28
rect 1369 22 1374 83
rect 1029 20 1034 21
rect 1028 19 1070 20
rect 1369 19 1372 22
rect 1384 19 1415 23
rect 1028 16 1372 19
rect 1028 13 1033 16
rect 1029 11 1033 13
rect 999 -11 1019 -7
rect 999 -20 1003 -11
rect 1021 -26 1023 -20
rect 1018 -67 1023 -26
rect 757 -106 765 -102
rect 770 -104 775 -102
rect 770 -106 997 -104
rect 365 -122 502 -117
rect 367 -123 376 -122
rect 577 -125 580 -117
rect 504 -128 515 -126
rect 577 -128 591 -125
rect 504 -129 509 -128
rect 285 -132 509 -129
rect 513 -132 515 -128
rect 285 -133 515 -132
rect 615 -134 618 -107
rect 677 -116 680 -106
rect 771 -107 997 -106
rect 784 -108 997 -107
rect 983 -116 987 -115
rect 677 -120 987 -116
rect 630 -128 689 -125
rect 520 -137 618 -134
rect 717 -128 979 -125
rect 703 -132 707 -129
rect 703 -135 770 -132
rect 208 -141 261 -140
rect 126 -144 261 -141
rect 520 -142 524 -137
rect 126 -150 129 -144
rect 75 -153 140 -150
rect 42 -169 83 -165
rect 79 -176 83 -169
rect 32 -208 33 -204
rect 40 -178 43 -177
rect 40 -181 47 -178
rect 40 -246 43 -181
rect 83 -180 116 -177
rect 136 -177 139 -153
rect 218 -153 303 -150
rect 307 -153 328 -150
rect 404 -151 469 -148
rect 272 -158 321 -157
rect 272 -160 317 -158
rect 272 -169 275 -160
rect 187 -181 220 -178
rect 200 -185 203 -181
rect 312 -185 315 -179
rect 200 -188 315 -185
rect 276 -197 277 -194
rect 274 -245 277 -197
rect 325 -203 328 -153
rect 465 -154 469 -151
rect 520 -154 523 -142
rect 766 -145 770 -135
rect 527 -148 547 -146
rect 527 -149 543 -148
rect 527 -153 528 -149
rect 532 -152 543 -149
rect 547 -151 632 -148
rect 731 -148 796 -145
rect 532 -153 547 -152
rect 527 -154 535 -153
rect 465 -157 523 -154
rect 369 -179 376 -176
rect 319 -207 353 -203
rect 313 -208 353 -207
rect 40 -249 134 -246
rect 144 -248 287 -245
rect 131 -253 134 -249
rect 303 -253 307 -221
rect 306 -256 307 -253
rect 282 -279 313 -275
rect 263 -280 287 -279
rect 220 -283 287 -280
rect 220 -284 223 -283
rect 164 -287 223 -284
rect 164 -296 168 -287
rect 74 -299 168 -296
rect 39 -327 46 -324
rect 39 -392 42 -327
rect 82 -326 115 -323
rect 135 -323 138 -299
rect 217 -299 302 -296
rect 271 -305 274 -303
rect 271 -308 318 -305
rect 96 -361 99 -326
rect 186 -327 219 -324
rect 199 -331 202 -327
rect 311 -331 314 -325
rect 199 -334 314 -331
rect 275 -343 276 -340
rect 196 -359 199 -343
rect 96 -365 189 -361
rect 195 -362 262 -359
rect 184 -378 189 -365
rect 184 -382 257 -378
rect 273 -391 276 -343
rect 326 -347 329 -208
rect 337 -231 358 -227
rect 369 -244 372 -179
rect 412 -178 445 -175
rect 465 -175 468 -157
rect 604 -159 762 -156
rect 688 -166 747 -163
rect 430 -227 434 -178
rect 516 -179 549 -176
rect 529 -183 532 -179
rect 641 -183 644 -177
rect 529 -186 644 -183
rect 688 -185 692 -166
rect 660 -189 692 -185
rect 696 -176 703 -173
rect 605 -195 606 -192
rect 443 -219 444 -216
rect 449 -219 540 -216
rect 603 -243 606 -195
rect 646 -205 680 -201
rect 640 -206 680 -205
rect 629 -223 633 -219
rect 369 -247 463 -244
rect 473 -246 606 -243
rect 630 -247 633 -223
rect 656 -234 684 -231
rect 696 -241 699 -176
rect 739 -175 772 -172
rect 792 -172 795 -148
rect 874 -148 959 -145
rect 851 -156 925 -154
rect 851 -157 929 -156
rect 745 -222 748 -191
rect 717 -225 748 -222
rect 755 -230 759 -175
rect 843 -176 876 -173
rect 856 -180 859 -176
rect 968 -180 971 -174
rect 856 -183 971 -180
rect 764 -217 767 -192
rect 932 -192 933 -189
rect 781 -229 840 -226
rect 848 -230 852 -192
rect 930 -240 933 -192
rect 696 -244 790 -241
rect 800 -243 943 -240
rect 460 -251 463 -247
rect 787 -248 790 -244
rect 337 -259 443 -255
rect 738 -255 742 -254
rect 677 -257 742 -255
rect 758 -255 778 -252
rect 758 -257 761 -255
rect 518 -258 761 -257
rect 518 -260 681 -258
rect 738 -260 761 -258
rect 775 -256 778 -255
rect 838 -255 886 -252
rect 775 -260 777 -256
rect 781 -260 782 -257
rect 518 -276 521 -260
rect 686 -266 687 -262
rect 691 -266 696 -263
rect 686 -267 696 -266
rect 700 -267 705 -263
rect 838 -264 841 -255
rect 769 -266 841 -264
rect 765 -267 841 -266
rect 847 -273 852 -270
rect 338 -279 521 -276
rect 547 -277 852 -273
rect 547 -278 670 -277
rect 548 -294 553 -278
rect 880 -291 883 -255
rect 964 -272 972 -269
rect 403 -297 468 -294
rect 337 -308 361 -305
rect 357 -328 361 -308
rect 435 -313 438 -297
rect 368 -325 375 -322
rect 357 -331 363 -328
rect 321 -348 351 -347
rect 321 -353 350 -348
rect 291 -382 311 -378
rect 39 -395 133 -392
rect 143 -394 286 -391
rect 130 -399 133 -395
rect 297 -406 312 -403
rect 322 -468 328 -353
rect 360 -369 363 -331
rect 349 -378 353 -377
rect 337 -382 353 -378
rect 333 -415 337 -406
rect 349 -403 353 -382
rect 368 -390 371 -325
rect 411 -324 444 -321
rect 464 -321 467 -297
rect 546 -297 631 -294
rect 730 -294 795 -291
rect 673 -302 751 -299
rect 674 -311 678 -302
rect 755 -302 757 -299
rect 604 -314 678 -311
rect 384 -377 388 -361
rect 411 -367 421 -365
rect 411 -369 416 -367
rect 415 -373 416 -369
rect 415 -374 421 -373
rect 426 -371 429 -324
rect 515 -325 548 -322
rect 528 -329 531 -325
rect 640 -329 643 -323
rect 528 -332 643 -329
rect 695 -322 702 -319
rect 435 -337 438 -336
rect 604 -341 605 -338
rect 435 -363 438 -341
rect 450 -359 588 -356
rect 426 -375 525 -371
rect 602 -389 605 -341
rect 644 -351 680 -348
rect 618 -375 677 -370
rect 695 -387 698 -322
rect 738 -321 771 -318
rect 791 -318 794 -294
rect 873 -294 958 -291
rect 968 -300 972 -272
rect 928 -303 972 -300
rect 928 -307 931 -303
rect 749 -348 753 -334
rect 722 -352 753 -348
rect 722 -362 726 -352
rect 749 -353 753 -352
rect 758 -357 762 -321
rect 842 -322 875 -319
rect 855 -326 858 -322
rect 967 -326 970 -320
rect 855 -329 970 -326
rect 931 -338 932 -335
rect 742 -361 762 -357
rect 758 -362 762 -361
rect 703 -366 726 -362
rect 703 -379 707 -366
rect 716 -373 843 -370
rect 849 -373 850 -370
rect 716 -374 850 -373
rect 703 -383 754 -379
rect 929 -386 932 -338
rect 950 -360 958 -358
rect 950 -364 952 -360
rect 957 -364 958 -360
rect 950 -366 958 -364
rect 368 -393 462 -390
rect 472 -392 615 -389
rect 669 -390 682 -388
rect 695 -390 789 -387
rect 799 -389 942 -386
rect 907 -390 920 -389
rect 459 -397 462 -393
rect 637 -391 682 -390
rect 637 -392 681 -391
rect 637 -394 674 -392
rect 678 -396 681 -392
rect 786 -394 789 -390
rect 678 -398 727 -396
rect 678 -400 719 -398
rect 349 -407 426 -403
rect 423 -411 426 -407
rect 506 -408 508 -403
rect 717 -404 719 -400
rect 724 -400 727 -398
rect 738 -398 742 -397
rect 724 -404 726 -400
rect 686 -408 687 -405
rect 717 -406 726 -404
rect 754 -402 757 -400
rect 506 -411 511 -408
rect 333 -416 385 -415
rect 333 -419 389 -416
rect 407 -440 411 -415
rect 423 -415 511 -411
rect 423 -416 426 -415
rect 686 -426 691 -408
rect 686 -429 723 -426
rect 688 -430 723 -429
rect 604 -431 609 -430
rect 738 -447 742 -402
rect 513 -450 742 -447
rect 513 -451 738 -450
rect 754 -452 757 -407
rect 907 -414 909 -408
rect 915 -414 916 -408
rect 907 -416 916 -414
rect 836 -451 843 -447
rect 950 -451 954 -366
rect 976 -408 979 -128
rect 836 -452 954 -451
rect 754 -455 954 -452
rect 975 -460 979 -408
rect 480 -464 514 -460
rect 569 -463 979 -460
rect 975 -464 979 -463
rect 510 -468 514 -464
rect 322 -496 325 -468
rect 510 -471 579 -468
rect 576 -475 579 -471
rect 983 -475 987 -120
rect 336 -480 379 -477
rect 384 -481 472 -477
rect 477 -481 557 -478
rect 576 -479 987 -475
rect 994 -489 997 -108
rect 1019 -141 1023 -67
rect 1029 -173 1034 11
rect 1131 10 1135 11
rect 1053 9 1262 10
rect 1425 9 1429 199
rect 1053 6 1429 9
rect 1109 -11 1112 -1
rect 1053 -36 1057 -18
rect 1053 -38 1099 -36
rect 1053 -39 1103 -38
rect 1109 -67 1112 -16
rect 1131 -20 1135 6
rect 1184 5 1429 6
rect 1312 4 1429 5
rect 1489 189 1511 193
rect 1300 -17 1301 -13
rect 1305 -17 1465 -13
rect 1185 -23 1194 -22
rect 1185 -26 1428 -23
rect 1131 -28 1135 -27
rect 1111 -87 1191 -84
rect 1111 -93 1114 -87
rect 403 -492 997 -489
rect 1002 -178 1034 -173
rect 1002 -391 1005 -178
rect 1019 -209 1023 -192
rect 1040 -194 1044 -95
rect 1072 -96 1114 -93
rect 1187 -94 1190 -87
rect 1211 -89 1270 -86
rect 1144 -97 1165 -94
rect 1191 -97 1217 -94
rect 1221 -97 1222 -94
rect 1267 -95 1270 -89
rect 1291 -94 1310 -91
rect 1267 -98 1274 -95
rect 1291 -99 1294 -94
rect 1314 -93 1353 -92
rect 1314 -95 1349 -93
rect 1087 -107 1099 -104
rect 1096 -171 1099 -107
rect 1159 -107 1241 -104
rect 1304 -104 1363 -101
rect 1274 -109 1277 -106
rect 1274 -112 1332 -109
rect 1423 -111 1426 -26
rect 1263 -131 1267 -113
rect 1423 -116 1446 -111
rect 1144 -135 1267 -131
rect 1144 -161 1148 -135
rect 1263 -136 1267 -135
rect 1412 -146 1447 -143
rect 1412 -147 1452 -146
rect 1278 -150 1336 -147
rect 1163 -155 1245 -152
rect 1278 -153 1281 -150
rect 1308 -158 1367 -155
rect 1148 -165 1169 -162
rect 1195 -165 1221 -162
rect 1225 -165 1226 -162
rect 1271 -164 1278 -161
rect 1191 -171 1194 -165
rect 1096 -174 1194 -171
rect 1271 -170 1274 -164
rect 1318 -166 1353 -164
rect 1460 -164 1465 -17
rect 1489 -141 1493 189
rect 1520 171 1523 218
rect 1527 218 1530 348
rect 1541 234 1545 396
rect 1595 383 1598 409
rect 1622 399 1625 417
rect 1553 380 1598 383
rect 1553 244 1556 380
rect 1595 376 1598 380
rect 1560 230 1563 367
rect 1622 356 1625 395
rect 1644 392 1647 494
rect 1782 486 1785 503
rect 1677 483 1785 486
rect 1644 389 1652 392
rect 1649 364 1652 389
rect 1598 353 1625 356
rect 1622 352 1625 353
rect 1632 361 1652 364
rect 1661 377 1664 462
rect 1677 433 1680 483
rect 1690 471 1699 474
rect 1661 364 1664 373
rect 1661 361 1680 364
rect 1632 345 1635 361
rect 1609 342 1635 345
rect 1639 354 1660 357
rect 1594 292 1597 305
rect 1609 293 1612 342
rect 1639 298 1642 354
rect 1677 349 1680 361
rect 1665 346 1680 349
rect 1689 362 1692 379
rect 1696 362 1699 471
rect 1756 436 1759 446
rect 1705 435 1759 436
rect 1708 433 1759 435
rect 1689 359 1699 362
rect 1689 346 1692 359
rect 1707 354 1725 357
rect 1665 314 1668 346
rect 1587 289 1597 292
rect 1527 216 1578 218
rect 1527 215 1581 216
rect 1560 195 1563 204
rect 1530 192 1563 195
rect 1518 168 1526 171
rect 1510 86 1514 143
rect 1523 132 1526 168
rect 1530 101 1533 192
rect 1587 180 1590 289
rect 1594 272 1597 289
rect 1604 290 1612 293
rect 1622 295 1642 298
rect 1653 311 1668 314
rect 1604 220 1607 290
rect 1622 278 1625 295
rect 1622 189 1625 274
rect 1653 188 1656 311
rect 1756 303 1759 433
rect 1661 298 1664 299
rect 1661 295 1688 298
rect 1661 255 1664 295
rect 1757 290 1764 293
rect 1688 257 1691 275
rect 1661 251 1672 255
rect 1661 234 1664 251
rect 1669 201 1672 251
rect 1688 254 1744 257
rect 1688 242 1691 254
rect 1689 202 1692 206
rect 1757 202 1760 290
rect 1795 276 1798 503
rect 1840 483 1844 531
rect 1830 478 1844 483
rect 1765 273 1798 276
rect 1765 229 1768 273
rect 1764 226 1769 229
rect 1669 198 1678 201
rect 1689 199 1760 202
rect 1653 184 1670 188
rect 1587 177 1596 180
rect 1666 165 1670 184
rect 1538 160 1670 165
rect 1538 105 1541 160
rect 1675 133 1678 198
rect 1690 191 1726 192
rect 1690 187 1717 191
rect 1690 144 1698 187
rect 1725 187 1726 191
rect 1766 161 1769 226
rect 1729 158 1769 161
rect 1774 152 1777 252
rect 1773 147 1826 152
rect 1697 138 1698 144
rect 1552 128 1635 132
rect 1675 130 1738 133
rect 1525 98 1533 101
rect 1506 82 1514 86
rect 1528 89 1599 92
rect 1489 -151 1493 -147
rect 1506 -150 1509 82
rect 1528 1 1531 89
rect 1596 85 1599 89
rect 1524 -2 1531 1
rect 1357 -166 1394 -164
rect 1318 -167 1394 -166
rect 1215 -173 1274 -170
rect 1040 -195 1233 -194
rect 1040 -196 1289 -195
rect 1040 -199 1376 -196
rect 1019 -212 1128 -209
rect 1019 -213 1023 -212
rect 1109 -232 1189 -229
rect 1109 -238 1112 -232
rect 1070 -241 1112 -238
rect 1185 -239 1188 -232
rect 1209 -234 1268 -231
rect 1142 -242 1163 -239
rect 1189 -242 1215 -239
rect 1219 -242 1220 -239
rect 1265 -240 1268 -234
rect 1289 -239 1308 -236
rect 1265 -243 1272 -240
rect 1289 -244 1292 -239
rect 1312 -238 1351 -237
rect 1312 -240 1347 -238
rect 1085 -252 1097 -249
rect 1094 -316 1097 -252
rect 1157 -252 1239 -249
rect 1302 -249 1361 -246
rect 1272 -254 1275 -251
rect 1272 -257 1330 -254
rect 1261 -276 1265 -258
rect 1373 -268 1376 -199
rect 1142 -280 1265 -276
rect 1142 -306 1146 -280
rect 1261 -281 1265 -280
rect 1322 -271 1376 -268
rect 1390 -267 1394 -167
rect 1460 -168 1472 -164
rect 1468 -252 1472 -168
rect 1505 -215 1509 -150
rect 1529 -142 1532 -12
rect 1538 -40 1541 75
rect 1579 65 1592 68
rect 1579 63 1582 65
rect 1556 60 1582 63
rect 1546 39 1580 43
rect 1546 -123 1550 39
rect 1589 32 1592 65
rect 1588 28 1592 32
rect 1597 23 1600 49
rect 1624 43 1627 57
rect 1611 39 1627 43
rect 1557 19 1600 23
rect 1557 -130 1561 19
rect 1597 16 1600 19
rect 1571 8 1574 11
rect 1606 8 1609 24
rect 1571 5 1609 8
rect 1571 -63 1574 5
rect 1624 -4 1627 39
rect 1600 -7 1627 -4
rect 1624 -8 1627 -7
rect 1632 -16 1635 128
rect 1735 127 1738 130
rect 1735 124 1813 127
rect 1679 121 1727 122
rect 1679 119 1724 121
rect 1663 17 1666 102
rect 1679 75 1682 119
rect 1692 111 1701 114
rect 1663 4 1666 13
rect 1663 1 1682 4
rect 1613 -19 1635 -16
rect 1641 -6 1662 -3
rect 1571 -64 1584 -63
rect 1571 -67 1581 -64
rect 1596 -68 1599 -55
rect 1589 -71 1599 -68
rect 1529 -144 1580 -142
rect 1529 -145 1583 -144
rect 1529 -155 1532 -145
rect 1589 -180 1592 -71
rect 1596 -88 1599 -71
rect 1606 -140 1609 -68
rect 1613 -78 1616 -19
rect 1641 -62 1644 -6
rect 1679 -11 1682 1
rect 1667 -14 1682 -11
rect 1691 2 1694 19
rect 1698 2 1701 111
rect 1758 76 1761 86
rect 1707 75 1761 76
rect 1710 73 1761 75
rect 1691 -1 1701 2
rect 1691 -14 1694 -1
rect 1709 -6 1727 -3
rect 1667 -46 1670 -14
rect 1624 -65 1644 -62
rect 1655 -49 1670 -46
rect 1613 -82 1617 -78
rect 1624 -82 1627 -65
rect 1589 -183 1598 -180
rect 1614 -196 1617 -82
rect 1624 -171 1627 -86
rect 1655 -172 1658 -49
rect 1758 -57 1761 73
rect 1663 -62 1666 -61
rect 1663 -65 1690 -62
rect 1663 -98 1666 -65
rect 1759 -70 1766 -67
rect 1663 -101 1680 -98
rect 1663 -126 1666 -101
rect 1655 -176 1672 -172
rect 1614 -199 1623 -196
rect 1499 -217 1509 -215
rect 1499 -223 1501 -217
rect 1507 -221 1509 -217
rect 1507 -223 1508 -221
rect 1499 -224 1508 -223
rect 1522 -236 1603 -231
rect 1471 -256 1472 -252
rect 1556 -259 1560 -250
rect 1556 -260 1557 -259
rect 1470 -261 1557 -260
rect 1469 -264 1557 -261
rect 1596 -261 1603 -236
rect 1620 -237 1623 -199
rect 1642 -229 1647 -186
rect 1668 -193 1672 -176
rect 1677 -227 1680 -101
rect 1690 -101 1693 -85
rect 1690 -104 1739 -101
rect 1690 -118 1693 -104
rect 1691 -158 1694 -154
rect 1759 -158 1762 -70
rect 1781 -106 1801 -102
rect 1777 -107 1801 -106
rect 1691 -161 1762 -158
rect 1692 -169 1728 -168
rect 1692 -173 1719 -169
rect 1692 -216 1700 -173
rect 1727 -173 1728 -169
rect 1722 -200 1753 -196
rect 1767 -197 1771 -153
rect 1699 -222 1700 -216
rect 1677 -230 1729 -227
rect 1620 -238 1638 -237
rect 1666 -238 1723 -235
rect 1620 -242 1670 -238
rect 1620 -261 1624 -260
rect 1390 -270 1401 -267
rect 1405 -270 1410 -267
rect 1322 -282 1325 -271
rect 1372 -278 1389 -275
rect 1386 -286 1389 -278
rect 1386 -290 1392 -286
rect 1396 -290 1397 -287
rect 1276 -295 1334 -292
rect 1161 -300 1243 -297
rect 1276 -298 1279 -295
rect 1306 -303 1365 -300
rect 1146 -310 1167 -307
rect 1193 -310 1219 -307
rect 1223 -310 1224 -307
rect 1269 -309 1276 -306
rect 1189 -316 1192 -310
rect 1094 -319 1192 -316
rect 1269 -315 1272 -309
rect 1316 -311 1351 -309
rect 1355 -311 1393 -309
rect 1316 -312 1393 -311
rect 1213 -318 1272 -315
rect 1312 -331 1376 -328
rect 1041 -332 1056 -331
rect 1046 -333 1056 -332
rect 1046 -334 1263 -333
rect 1312 -334 1315 -331
rect 1046 -336 1315 -334
rect 1041 -337 1315 -336
rect 1020 -352 1024 -351
rect 1020 -355 1127 -352
rect 1020 -391 1024 -355
rect 1322 -366 1325 -339
rect 1110 -374 1190 -371
rect 1110 -380 1113 -374
rect 1071 -383 1113 -380
rect 1186 -381 1189 -374
rect 1210 -376 1269 -373
rect 1125 -385 1139 -382
rect 1143 -384 1164 -381
rect 1143 -385 1145 -384
rect 1190 -384 1216 -381
rect 1220 -384 1221 -381
rect 1266 -382 1269 -376
rect 1290 -381 1309 -378
rect 1266 -385 1273 -382
rect 1002 -394 1026 -391
rect 1086 -394 1098 -391
rect 1002 -453 1005 -394
rect 1071 -431 1073 -427
rect 1002 -456 1009 -453
rect 1068 -453 1072 -431
rect 1013 -456 1072 -453
rect 1002 -493 1005 -456
rect 1095 -458 1098 -394
rect 1125 -396 1128 -385
rect 1290 -386 1293 -381
rect 1313 -380 1352 -379
rect 1313 -382 1348 -380
rect 1158 -394 1240 -391
rect 1303 -391 1362 -388
rect 1273 -396 1276 -393
rect 1106 -399 1128 -396
rect 1106 -426 1109 -399
rect 1273 -399 1331 -396
rect 1262 -418 1266 -400
rect 1373 -403 1376 -331
rect 1390 -357 1393 -312
rect 1390 -360 1404 -357
rect 1408 -360 1413 -357
rect 1469 -403 1472 -264
rect 1556 -265 1560 -264
rect 1596 -268 1624 -261
rect 1322 -409 1323 -405
rect 1373 -406 1473 -403
rect 1373 -409 1376 -406
rect 1143 -422 1266 -418
rect 1143 -448 1147 -422
rect 1262 -423 1266 -422
rect 1320 -422 1323 -409
rect 1501 -410 1506 -283
rect 1408 -418 1411 -411
rect 1373 -421 1411 -418
rect 1320 -424 1325 -422
rect 1320 -426 1321 -424
rect 1277 -437 1335 -434
rect 1162 -442 1244 -439
rect 1277 -440 1280 -437
rect 1307 -445 1366 -442
rect 1391 -445 1397 -442
rect 1401 -445 1414 -442
rect 1147 -452 1168 -449
rect 1194 -452 1220 -449
rect 1224 -452 1225 -449
rect 1270 -451 1277 -448
rect 1190 -458 1193 -452
rect 1095 -461 1193 -458
rect 1270 -457 1273 -451
rect 1317 -453 1352 -451
rect 1317 -454 1356 -453
rect 1214 -460 1273 -457
rect 1345 -458 1348 -454
rect 1391 -458 1394 -445
rect 1345 -461 1394 -458
rect 1321 -483 1322 -479
rect 1055 -489 1059 -488
rect 322 -503 323 -496
rect 625 -501 626 -497
rect 630 -499 633 -497
rect 630 -501 1004 -499
rect 625 -502 1004 -501
rect 907 -538 911 -532
rect 916 -538 940 -532
rect 907 -540 940 -538
rect 996 -548 999 -502
rect 1055 -523 1059 -494
rect 1054 -524 1195 -523
rect 1054 -528 1306 -524
rect 995 -555 1013 -548
rect 996 -557 999 -555
rect 1321 -562 1324 -483
rect 1321 -566 1355 -562
rect 1360 -566 1367 -562
rect 1454 -576 1460 -478
rect 1501 -536 1504 -410
rect 1587 -498 1593 -496
rect 1590 -505 1593 -498
rect 1587 -535 1593 -505
rect 1607 -522 1611 -507
rect 1491 -541 1504 -536
rect 1582 -539 1594 -535
rect 1582 -545 1584 -539
rect 1590 -545 1594 -539
rect 1582 -547 1594 -545
rect 1620 -551 1624 -268
rect 1655 -339 1658 -254
rect 1666 -281 1670 -242
rect 1684 -245 1693 -242
rect 1666 -284 1667 -281
rect 1683 -354 1686 -337
rect 1690 -354 1693 -245
rect 1720 -273 1723 -238
rect 1750 -262 1753 -200
rect 1783 -227 1787 -226
rect 1762 -230 1787 -227
rect 1734 -266 1753 -262
rect 1720 -276 1775 -273
rect 1699 -281 1753 -280
rect 1702 -283 1753 -281
rect 1737 -303 1740 -295
rect 1726 -306 1740 -303
rect 1726 -334 1729 -306
rect 1683 -357 1693 -354
rect 1683 -370 1686 -357
rect 1702 -364 1729 -360
rect 1655 -418 1658 -417
rect 1655 -421 1682 -418
rect 1655 -482 1658 -421
rect 1700 -429 1704 -364
rect 1711 -371 1714 -368
rect 1711 -374 1718 -371
rect 1711 -422 1714 -374
rect 1726 -378 1729 -364
rect 1725 -381 1729 -378
rect 1725 -417 1728 -381
rect 1750 -406 1753 -283
rect 1747 -409 1753 -406
rect 1747 -410 1750 -409
rect 1733 -413 1750 -410
rect 1758 -417 1776 -413
rect 1711 -425 1721 -422
rect 1736 -424 1743 -421
rect 1700 -432 1732 -429
rect 1700 -433 1728 -432
rect 1682 -457 1685 -441
rect 1662 -460 1685 -457
rect 1635 -507 1636 -503
rect 1633 -528 1636 -507
rect 1633 -532 1653 -528
rect 1620 -554 1654 -551
rect 1582 -558 1602 -554
rect 1480 -566 1640 -562
rect 1663 -572 1666 -460
rect 1682 -474 1685 -460
rect 1701 -492 1704 -449
rect 1675 -495 1704 -492
rect 1675 -550 1678 -495
rect 1725 -497 1728 -433
rect 1736 -468 1739 -424
rect 1773 -426 1776 -417
rect 1751 -429 1776 -426
rect 1736 -472 1740 -468
rect 1683 -514 1686 -510
rect 1751 -514 1754 -429
rect 1683 -517 1754 -514
rect 1693 -547 1697 -532
rect 1766 -550 1769 -443
rect 1675 -570 1678 -555
rect 1716 -557 1718 -553
rect 1722 -557 1729 -553
rect 1716 -558 1729 -557
rect 1759 -553 1769 -550
rect 1716 -560 1732 -558
rect 1766 -564 1769 -553
rect 1453 -577 1474 -576
rect 1453 -579 1617 -577
rect 1783 -579 1787 -230
rect 1795 -562 1801 -107
rect 1808 -313 1813 124
rect 1820 -36 1826 147
rect 1820 -102 1827 -36
rect 1800 -566 1801 -562
rect 1807 -574 1813 -313
rect 1821 -563 1827 -102
rect 1831 -304 1835 478
rect 1821 -565 1832 -563
rect 1821 -571 1823 -565
rect 1830 -571 1832 -565
rect 1821 -572 1832 -571
rect 1453 -580 1657 -579
rect 1673 -580 1789 -579
rect 1453 -581 1789 -580
rect 1611 -583 1789 -581
<< metal3 >>
rect 497 378 522 380
rect 497 374 498 378
rect 502 374 522 378
rect 497 373 503 374
rect 516 359 522 374
rect 516 357 523 359
rect 516 353 517 357
rect 521 353 523 357
rect 516 352 523 353
rect 1433 308 1491 309
rect 1433 303 1435 308
rect 1440 303 1491 308
rect 1433 302 1491 303
rect 1484 286 1491 302
rect 1484 285 1522 286
rect 1484 280 1515 285
rect 1520 280 1522 285
rect 1514 279 1522 280
rect 1299 43 1306 44
rect 1299 38 1300 43
rect 1305 38 1306 43
rect 1299 37 1306 38
rect 1013 33 1020 34
rect 1013 28 1014 33
rect 1019 28 1020 33
rect 278 13 293 14
rect -43 12 293 13
rect -43 7 283 12
rect -42 -104 -36 7
rect 278 5 283 7
rect 289 5 293 12
rect 278 2 293 5
rect 1013 3 1020 28
rect 1013 -3 1188 3
rect 1180 -14 1186 -3
rect 1178 -19 1186 -14
rect 1300 -13 1306 37
rect 1300 -17 1301 -13
rect 1305 -17 1306 -13
rect 1300 -18 1306 -17
rect 1178 -26 1179 -19
rect 1185 -26 1186 -19
rect 1178 -27 1186 -26
rect -15 -104 -6 -102
rect -42 -105 -6 -104
rect -42 -110 -12 -105
rect -8 -110 -6 -105
rect -15 -113 -6 -110
rect 521 -104 531 -103
rect 521 -108 525 -104
rect 529 -108 531 -104
rect 521 -109 531 -108
rect 521 -115 527 -109
rect 521 -121 661 -115
rect 508 -128 533 -126
rect 508 -132 509 -128
rect 513 -132 533 -128
rect 508 -133 514 -132
rect 527 -147 533 -132
rect 527 -149 534 -147
rect 527 -153 528 -149
rect 532 -153 534 -149
rect 527 -154 534 -153
rect 655 -184 661 -121
rect 655 -189 656 -184
rect 660 -189 661 -184
rect 655 -191 661 -189
rect 1499 -217 1508 -215
rect 1499 -223 1501 -217
rect 1507 -223 1508 -217
rect 1499 -224 1508 -223
rect 686 -262 692 -261
rect 686 -266 687 -262
rect 691 -266 692 -262
rect 686 -320 692 -266
rect 1500 -277 1507 -224
rect 1500 -283 1501 -277
rect 1506 -283 1507 -277
rect 1500 -285 1507 -283
rect 411 -367 422 -365
rect 411 -373 416 -367
rect 421 -373 422 -367
rect 411 -374 422 -373
rect 415 -425 422 -374
rect 685 -376 692 -320
rect 1005 -332 1047 -331
rect 1005 -336 1041 -332
rect 1046 -336 1047 -332
rect 1005 -337 1047 -336
rect 1005 -358 1011 -337
rect 950 -360 1011 -358
rect 950 -364 952 -360
rect 957 -364 1011 -360
rect 950 -366 1011 -364
rect 685 -401 691 -376
rect 717 -398 726 -396
rect 685 -404 697 -401
rect 685 -408 687 -404
rect 691 -408 697 -404
rect 717 -404 719 -398
rect 724 -400 726 -398
rect 913 -399 924 -395
rect 863 -400 924 -399
rect 724 -401 924 -400
rect 724 -403 922 -401
rect 724 -404 919 -403
rect 717 -407 919 -404
rect 685 -409 697 -408
rect 907 -408 918 -407
rect 907 -414 909 -408
rect 915 -414 918 -408
rect 907 -416 918 -414
rect 415 -426 633 -425
rect 415 -430 604 -426
rect 609 -430 633 -426
rect 415 -431 633 -430
rect 625 -497 633 -431
rect 625 -501 626 -497
rect 630 -501 633 -497
rect 625 -502 633 -501
rect 908 -532 918 -416
rect 908 -538 911 -532
rect 916 -538 918 -532
rect 908 -540 918 -538
rect 1582 -539 1723 -535
rect 1582 -545 1584 -539
rect 1590 -541 1723 -539
rect 1590 -545 1594 -541
rect 1582 -547 1594 -545
rect 1717 -553 1723 -541
rect 1600 -554 1607 -553
rect 1600 -558 1602 -554
rect 1606 -558 1607 -554
rect 1600 -567 1607 -558
rect 1717 -557 1718 -553
rect 1722 -557 1723 -553
rect 1717 -559 1723 -557
rect 1821 -565 1832 -563
rect 1821 -567 1823 -565
rect 1600 -571 1823 -567
rect 1830 -571 1832 -565
rect 1600 -573 1832 -571
rect 1821 -574 1832 -573
<< ntransistor >>
rect 1701 464 1710 466
rect 1701 457 1710 459
rect 121 425 123 436
rect 128 425 130 436
rect 141 425 143 434
rect 208 425 210 436
rect 215 425 217 436
rect 228 425 230 434
rect 301 425 303 436
rect 308 425 310 436
rect 321 425 323 434
rect 541 427 543 436
rect 554 427 556 438
rect 561 427 563 438
rect 634 427 636 436
rect 647 427 649 438
rect 654 427 656 438
rect 721 427 723 436
rect 734 427 736 438
rect 741 427 743 438
rect 1698 445 1704 447
rect 1582 436 1588 438
rect 1576 424 1585 426
rect 1576 417 1585 419
rect 1042 392 1044 395
rect 1698 418 1710 420
rect 1698 411 1710 413
rect 1698 401 1707 403
rect 1114 391 1116 394
rect 1153 391 1155 397
rect 1174 391 1176 397
rect 1207 391 1209 397
rect 1228 391 1230 397
rect 1263 391 1265 397
rect 1284 391 1286 397
rect 1317 391 1319 397
rect 1338 391 1340 397
rect 1698 391 1707 393
rect 1693 375 1702 377
rect 43 313 45 319
rect 55 307 57 316
rect 62 307 64 316
rect 121 315 123 324
rect 137 310 139 319
rect 147 310 149 319
rect 157 307 159 319
rect 164 307 166 319
rect 205 315 207 324
rect 221 310 223 319
rect 231 310 233 319
rect 241 307 243 319
rect 248 307 250 319
rect 275 313 277 319
rect 287 307 289 316
rect 294 307 296 316
rect 372 315 374 321
rect 384 309 386 318
rect 391 309 393 318
rect 450 317 452 326
rect 466 312 468 321
rect 476 312 478 321
rect 486 309 488 321
rect 493 309 495 321
rect 534 317 536 326
rect 550 312 552 321
rect 560 312 562 321
rect 570 309 572 321
rect 577 309 579 321
rect 604 315 606 321
rect 699 318 701 324
rect 1118 369 1120 372
rect 1157 366 1159 372
rect 1178 366 1180 372
rect 1211 366 1213 372
rect 1232 366 1234 372
rect 1267 366 1269 372
rect 1288 366 1290 372
rect 1321 366 1323 372
rect 1342 366 1344 372
rect 1584 358 1593 360
rect 616 309 618 318
rect 623 309 625 318
rect 711 312 713 321
rect 718 312 720 321
rect 777 320 779 329
rect 793 315 795 324
rect 803 315 805 324
rect 813 312 815 324
rect 820 312 822 324
rect 861 320 863 329
rect 877 315 879 324
rect 887 315 889 324
rect 897 312 899 324
rect 904 312 906 324
rect 931 318 933 324
rect 1548 343 1554 345
rect 1548 333 1554 335
rect 1548 323 1554 325
rect 943 312 945 321
rect 950 312 952 321
rect 1579 342 1588 344
rect 1579 332 1588 334
rect 1698 334 1710 336
rect 1698 327 1710 329
rect 1576 322 1588 324
rect 1576 315 1588 317
rect 1698 317 1707 319
rect 1698 307 1707 309
rect 136 279 138 285
rect 146 279 148 285
rect 156 279 158 285
rect 465 281 467 287
rect 475 281 477 287
rect 485 281 487 287
rect 792 284 794 290
rect 802 284 804 290
rect 812 284 814 290
rect 1732 326 1738 328
rect 1732 316 1738 318
rect 1732 306 1738 308
rect 1693 291 1702 293
rect 1584 274 1593 276
rect 1042 247 1044 250
rect 1383 254 1385 264
rect 1114 246 1116 249
rect 1153 246 1155 252
rect 1174 246 1176 252
rect 1207 246 1209 252
rect 1228 246 1230 252
rect 1263 246 1265 252
rect 1284 246 1286 252
rect 1317 246 1319 252
rect 1338 246 1340 252
rect 1395 250 1397 264
rect 1579 258 1588 260
rect 1579 248 1588 250
rect 1576 238 1588 240
rect 42 167 44 173
rect 54 161 56 170
rect 61 161 63 170
rect 120 169 122 178
rect 136 164 138 173
rect 146 164 148 173
rect 156 161 158 173
rect 163 161 165 173
rect 204 169 206 178
rect 220 164 222 173
rect 230 164 232 173
rect 240 161 242 173
rect 247 161 249 173
rect 274 167 276 173
rect 286 161 288 170
rect 293 161 295 170
rect 371 169 373 175
rect 383 163 385 172
rect 390 163 392 172
rect 449 171 451 180
rect 465 166 467 175
rect 475 166 477 175
rect 485 163 487 175
rect 492 163 494 175
rect 533 171 535 180
rect 549 166 551 175
rect 559 166 561 175
rect 569 163 571 175
rect 576 163 578 175
rect 603 169 605 175
rect 698 172 700 178
rect 1118 224 1120 227
rect 1157 221 1159 227
rect 1178 221 1180 227
rect 1211 221 1213 227
rect 1232 221 1234 227
rect 1267 221 1269 227
rect 1288 221 1290 227
rect 1321 221 1323 227
rect 1342 221 1344 227
rect 1576 231 1588 233
rect 1384 215 1386 225
rect 1396 215 1398 229
rect 1701 232 1710 234
rect 1701 225 1710 227
rect 1698 213 1704 215
rect 1582 204 1588 206
rect 615 163 617 172
rect 622 163 624 172
rect 710 166 712 175
rect 717 166 719 175
rect 776 174 778 183
rect 792 169 794 178
rect 802 169 804 178
rect 812 166 814 178
rect 819 166 821 178
rect 860 174 862 183
rect 876 169 878 178
rect 886 169 888 178
rect 896 166 898 178
rect 903 166 905 178
rect 930 172 932 178
rect 942 166 944 175
rect 949 166 951 175
rect 1576 192 1585 194
rect 1576 185 1585 187
rect 135 133 137 139
rect 145 133 147 139
rect 155 133 157 139
rect 464 135 466 141
rect 474 135 476 141
rect 484 135 486 141
rect 791 138 793 144
rect 801 138 803 144
rect 811 138 813 144
rect 1041 105 1043 108
rect 1383 114 1385 124
rect 1113 104 1115 107
rect 1152 104 1154 110
rect 1173 104 1175 110
rect 1206 104 1208 110
rect 1227 104 1229 110
rect 1262 104 1264 110
rect 1283 104 1285 110
rect 1316 104 1318 110
rect 1337 104 1339 110
rect 1395 110 1397 124
rect 1703 104 1712 106
rect 1703 97 1712 99
rect 1117 82 1119 85
rect 1156 79 1158 85
rect 1177 79 1179 85
rect 1210 79 1212 85
rect 1231 79 1233 85
rect 1266 79 1268 85
rect 1287 79 1289 85
rect 1320 79 1322 85
rect 1341 79 1343 85
rect 1700 85 1706 87
rect 1584 76 1590 78
rect 1578 64 1587 66
rect 1578 57 1587 59
rect 1700 58 1712 60
rect 1700 51 1712 53
rect 1700 41 1709 43
rect 1700 31 1709 33
rect 336 19 338 28
rect 349 17 351 28
rect 356 17 358 28
rect 429 19 431 28
rect 442 17 444 28
rect 449 17 451 28
rect 516 19 518 28
rect 529 17 531 28
rect 536 17 538 28
rect 1695 15 1704 17
rect 1586 -2 1595 0
rect 1550 -17 1556 -15
rect 1550 -27 1556 -25
rect 1550 -37 1556 -35
rect 1581 -18 1590 -16
rect 1581 -28 1590 -26
rect 1700 -26 1712 -24
rect 1700 -33 1712 -31
rect 1578 -38 1590 -36
rect 1578 -45 1590 -43
rect 1700 -43 1709 -41
rect 1700 -53 1709 -51
rect 132 -81 134 -70
rect 139 -81 141 -70
rect 152 -81 154 -72
rect 219 -81 221 -70
rect 226 -81 228 -70
rect 239 -81 241 -72
rect 312 -81 314 -70
rect 319 -81 321 -70
rect 332 -81 334 -72
rect 552 -79 554 -70
rect 565 -79 567 -68
rect 572 -79 574 -68
rect 645 -79 647 -70
rect 658 -79 660 -68
rect 665 -79 667 -68
rect 1734 -34 1740 -32
rect 1734 -44 1740 -42
rect 1734 -54 1740 -52
rect 732 -79 734 -70
rect 745 -79 747 -68
rect 752 -79 754 -68
rect 1695 -69 1704 -67
rect 1586 -86 1595 -84
rect 1063 -119 1065 -116
rect 1581 -102 1590 -100
rect 1581 -112 1590 -110
rect 1135 -120 1137 -117
rect 1174 -120 1176 -114
rect 1195 -120 1197 -114
rect 1228 -120 1230 -114
rect 1249 -120 1251 -114
rect 1284 -120 1286 -114
rect 1305 -120 1307 -114
rect 1338 -120 1340 -114
rect 1359 -120 1361 -114
rect 1578 -122 1590 -120
rect 1578 -129 1590 -127
rect 54 -193 56 -187
rect 66 -199 68 -190
rect 73 -199 75 -190
rect 132 -191 134 -182
rect 148 -196 150 -187
rect 158 -196 160 -187
rect 168 -199 170 -187
rect 175 -199 177 -187
rect 216 -191 218 -182
rect 232 -196 234 -187
rect 242 -196 244 -187
rect 252 -199 254 -187
rect 259 -199 261 -187
rect 286 -193 288 -187
rect 298 -199 300 -190
rect 305 -199 307 -190
rect 383 -191 385 -185
rect 395 -197 397 -188
rect 402 -197 404 -188
rect 461 -189 463 -180
rect 477 -194 479 -185
rect 487 -194 489 -185
rect 497 -197 499 -185
rect 504 -197 506 -185
rect 545 -189 547 -180
rect 561 -194 563 -185
rect 571 -194 573 -185
rect 581 -197 583 -185
rect 588 -197 590 -185
rect 615 -191 617 -185
rect 710 -188 712 -182
rect 1703 -128 1712 -126
rect 1703 -135 1712 -133
rect 1139 -142 1141 -139
rect 1178 -145 1180 -139
rect 1199 -145 1201 -139
rect 1232 -145 1234 -139
rect 1253 -145 1255 -139
rect 1288 -145 1290 -139
rect 1309 -145 1311 -139
rect 1342 -145 1344 -139
rect 1363 -145 1365 -139
rect 1700 -147 1706 -145
rect 1584 -156 1590 -154
rect 627 -197 629 -188
rect 634 -197 636 -188
rect 722 -194 724 -185
rect 729 -194 731 -185
rect 788 -186 790 -177
rect 804 -191 806 -182
rect 814 -191 816 -182
rect 824 -194 826 -182
rect 831 -194 833 -182
rect 872 -186 874 -177
rect 888 -191 890 -182
rect 898 -191 900 -182
rect 908 -194 910 -182
rect 915 -194 917 -182
rect 942 -188 944 -182
rect 1578 -168 1587 -166
rect 1578 -175 1587 -173
rect 954 -194 956 -185
rect 961 -194 963 -185
rect 147 -227 149 -221
rect 157 -227 159 -221
rect 167 -227 169 -221
rect 476 -225 478 -219
rect 486 -225 488 -219
rect 496 -225 498 -219
rect 803 -222 805 -216
rect 813 -222 815 -216
rect 823 -222 825 -216
rect 1061 -264 1063 -261
rect 1415 -258 1417 -248
rect 1427 -258 1429 -244
rect 1695 -252 1704 -250
rect 1133 -265 1135 -262
rect 1172 -265 1174 -259
rect 1193 -265 1195 -259
rect 1226 -265 1228 -259
rect 1247 -265 1249 -259
rect 1282 -265 1284 -259
rect 1303 -265 1305 -259
rect 1336 -265 1338 -259
rect 1357 -265 1359 -259
rect 1695 -259 1704 -257
rect 53 -339 55 -333
rect 65 -345 67 -336
rect 72 -345 74 -336
rect 131 -337 133 -328
rect 147 -342 149 -333
rect 157 -342 159 -333
rect 167 -345 169 -333
rect 174 -345 176 -333
rect 215 -337 217 -328
rect 231 -342 233 -333
rect 241 -342 243 -333
rect 251 -345 253 -333
rect 258 -345 260 -333
rect 285 -339 287 -333
rect 297 -345 299 -336
rect 304 -345 306 -336
rect 382 -337 384 -331
rect 394 -343 396 -334
rect 401 -343 403 -334
rect 460 -335 462 -326
rect 476 -340 478 -331
rect 486 -340 488 -331
rect 496 -343 498 -331
rect 503 -343 505 -331
rect 544 -335 546 -326
rect 560 -340 562 -331
rect 570 -340 572 -331
rect 580 -343 582 -331
rect 587 -343 589 -331
rect 614 -337 616 -331
rect 709 -334 711 -328
rect 1137 -287 1139 -284
rect 1176 -290 1178 -284
rect 1197 -290 1199 -284
rect 1230 -290 1232 -284
rect 1251 -290 1253 -284
rect 1286 -290 1288 -284
rect 1307 -290 1309 -284
rect 1340 -290 1342 -284
rect 1361 -290 1363 -284
rect 1692 -271 1698 -269
rect 1692 -298 1704 -296
rect 1692 -305 1704 -303
rect 626 -343 628 -334
rect 633 -343 635 -334
rect 721 -340 723 -331
rect 728 -340 730 -331
rect 787 -332 789 -323
rect 803 -337 805 -328
rect 813 -337 815 -328
rect 823 -340 825 -328
rect 830 -340 832 -328
rect 871 -332 873 -323
rect 887 -337 889 -328
rect 897 -337 899 -328
rect 907 -340 909 -328
rect 914 -340 916 -328
rect 941 -334 943 -328
rect 1692 -315 1701 -313
rect 1692 -325 1701 -323
rect 953 -340 955 -331
rect 960 -340 962 -331
rect 146 -373 148 -367
rect 156 -373 158 -367
rect 166 -373 168 -367
rect 475 -371 477 -365
rect 485 -371 487 -365
rect 495 -371 497 -365
rect 802 -368 804 -362
rect 812 -368 814 -362
rect 822 -368 824 -362
rect 1687 -341 1696 -339
rect 1417 -381 1419 -371
rect 1429 -385 1431 -371
rect 1062 -406 1064 -403
rect 1692 -382 1704 -380
rect 1692 -389 1704 -387
rect 1692 -399 1701 -397
rect 1134 -407 1136 -404
rect 1173 -407 1175 -401
rect 1194 -407 1196 -401
rect 1227 -407 1229 -401
rect 1248 -407 1250 -401
rect 1283 -407 1285 -401
rect 1304 -407 1306 -401
rect 1337 -407 1339 -401
rect 1358 -407 1360 -401
rect 1692 -409 1701 -407
rect 1138 -429 1140 -426
rect 1177 -432 1179 -426
rect 1198 -432 1200 -426
rect 1231 -432 1233 -426
rect 1252 -432 1254 -426
rect 1287 -432 1289 -426
rect 1308 -432 1310 -426
rect 1341 -432 1343 -426
rect 1362 -432 1364 -426
rect 1419 -437 1421 -427
rect 1431 -437 1433 -423
rect 1726 -390 1732 -388
rect 1726 -400 1732 -398
rect 1726 -410 1732 -408
rect 1687 -425 1696 -423
rect 1716 -438 1729 -436
rect 1719 -448 1729 -446
rect 347 -487 349 -478
rect 360 -489 362 -478
rect 367 -489 369 -478
rect 440 -487 442 -478
rect 453 -489 455 -478
rect 460 -489 462 -478
rect 527 -487 529 -478
rect 540 -489 542 -478
rect 547 -489 549 -478
rect 1722 -458 1736 -456
rect 1722 -468 1736 -466
rect 1695 -484 1704 -482
rect 1716 -488 1736 -486
rect 1695 -491 1704 -489
rect 1716 -495 1736 -493
rect 1692 -503 1698 -501
rect 1716 -506 1730 -504
<< ptransistor >>
rect 1671 465 1681 467
rect 1671 455 1681 457
rect 1042 428 1044 434
rect 1669 445 1681 447
rect 1114 428 1116 434
rect 1153 428 1155 434
rect 1174 428 1176 434
rect 1207 428 1209 434
rect 1228 428 1230 434
rect 1263 428 1265 434
rect 1284 428 1286 434
rect 1317 428 1319 434
rect 1338 428 1340 434
rect 1605 436 1617 438
rect 121 390 123 403
rect 131 390 133 403
rect 141 392 143 410
rect 208 390 210 403
rect 218 390 220 403
rect 228 392 230 410
rect 301 390 303 403
rect 311 390 313 403
rect 321 392 323 410
rect 541 394 543 412
rect 551 392 553 405
rect 561 392 563 405
rect 634 394 636 412
rect 644 392 646 405
rect 654 392 656 405
rect 721 394 723 412
rect 1605 426 1615 428
rect 731 392 733 405
rect 741 392 743 405
rect 1605 416 1615 418
rect 1653 419 1680 421
rect 1662 409 1680 411
rect 1662 399 1680 401
rect 1653 383 1680 385
rect 43 336 45 348
rect 53 336 55 346
rect 63 336 65 346
rect 129 337 131 364
rect 145 337 147 355
rect 155 337 157 355
rect 165 337 167 364
rect 213 337 215 364
rect 229 337 231 355
rect 239 337 241 355
rect 249 337 251 364
rect 275 336 277 348
rect 285 336 287 346
rect 295 336 297 346
rect 372 338 374 350
rect 382 338 384 348
rect 392 338 394 348
rect 458 339 460 366
rect 474 339 476 357
rect 484 339 486 357
rect 494 339 496 366
rect 542 339 544 366
rect 558 339 560 357
rect 568 339 570 357
rect 578 339 580 366
rect 604 338 606 350
rect 614 338 616 348
rect 624 338 626 348
rect 699 341 701 353
rect 709 341 711 351
rect 719 341 721 351
rect 785 342 787 369
rect 801 342 803 360
rect 811 342 813 360
rect 821 342 823 369
rect 869 342 871 369
rect 885 342 887 360
rect 895 342 897 360
rect 905 342 907 369
rect 931 341 933 353
rect 941 341 943 351
rect 951 341 953 351
rect 1503 343 1521 345
rect 1503 336 1521 338
rect 1118 329 1120 335
rect 1157 329 1159 335
rect 1178 329 1180 335
rect 1211 329 1213 335
rect 1232 329 1234 335
rect 1267 329 1269 335
rect 1288 329 1290 335
rect 1321 329 1323 335
rect 1342 329 1344 335
rect 1512 323 1524 325
rect 1606 350 1633 352
rect 1606 334 1624 336
rect 1653 335 1680 337
rect 1606 324 1624 326
rect 1662 325 1680 327
rect 1606 314 1633 316
rect 1662 315 1680 317
rect 136 234 138 252
rect 143 234 145 252
rect 156 243 158 255
rect 1042 283 1044 289
rect 1114 283 1116 289
rect 1153 283 1155 289
rect 1174 283 1176 289
rect 1207 283 1209 289
rect 1228 283 1230 289
rect 1263 283 1265 289
rect 1284 283 1286 289
rect 1317 283 1319 289
rect 1338 283 1340 289
rect 1383 276 1385 293
rect 1395 276 1397 304
rect 1653 299 1680 301
rect 1762 326 1774 328
rect 1765 313 1783 315
rect 1765 306 1783 308
rect 465 236 467 254
rect 472 236 474 254
rect 485 245 487 257
rect 792 239 794 257
rect 799 239 801 257
rect 812 248 814 260
rect 1606 266 1633 268
rect 1606 250 1624 252
rect 1606 240 1624 242
rect 42 190 44 202
rect 52 190 54 200
rect 62 190 64 200
rect 128 191 130 218
rect 144 191 146 209
rect 154 191 156 209
rect 164 191 166 218
rect 212 191 214 218
rect 228 191 230 209
rect 238 191 240 209
rect 248 191 250 218
rect 274 190 276 202
rect 284 190 286 200
rect 294 190 296 200
rect 371 192 373 204
rect 381 192 383 202
rect 391 192 393 202
rect 457 193 459 220
rect 473 193 475 211
rect 483 193 485 211
rect 493 193 495 220
rect 541 193 543 220
rect 557 193 559 211
rect 567 193 569 211
rect 577 193 579 220
rect 603 192 605 204
rect 613 192 615 202
rect 623 192 625 202
rect 698 195 700 207
rect 708 195 710 205
rect 718 195 720 205
rect 784 196 786 223
rect 800 196 802 214
rect 810 196 812 214
rect 820 196 822 223
rect 868 196 870 223
rect 884 196 886 214
rect 894 196 896 214
rect 904 196 906 223
rect 930 195 932 207
rect 1606 230 1633 232
rect 1671 233 1681 235
rect 1671 223 1681 225
rect 1669 213 1681 215
rect 940 195 942 205
rect 950 195 952 205
rect 1118 184 1120 190
rect 1157 184 1159 190
rect 1178 184 1180 190
rect 1211 184 1213 190
rect 1232 184 1234 190
rect 1267 184 1269 190
rect 1288 184 1290 190
rect 1321 184 1323 190
rect 1342 184 1344 190
rect 1384 186 1386 203
rect 1396 175 1398 203
rect 1605 204 1617 206
rect 1605 194 1615 196
rect 1605 184 1615 186
rect 1041 141 1043 147
rect 1113 141 1115 147
rect 1152 141 1154 147
rect 1173 141 1175 147
rect 1206 141 1208 147
rect 1227 141 1229 147
rect 1262 141 1264 147
rect 1283 141 1285 147
rect 1316 141 1318 147
rect 1337 141 1339 147
rect 135 88 137 106
rect 142 88 144 106
rect 155 97 157 109
rect 1383 136 1385 153
rect 1395 136 1397 164
rect 464 90 466 108
rect 471 90 473 108
rect 484 99 486 111
rect 791 93 793 111
rect 798 93 800 111
rect 811 102 813 114
rect 1673 105 1683 107
rect 1673 95 1683 97
rect 336 43 338 61
rect 346 50 348 63
rect 356 50 358 63
rect 429 43 431 61
rect 439 50 441 63
rect 449 50 451 63
rect 1671 85 1683 87
rect 1607 76 1619 78
rect 1607 66 1617 68
rect 516 43 518 61
rect 526 50 528 63
rect 536 50 538 63
rect 1607 56 1617 58
rect 1655 59 1682 61
rect 1664 49 1682 51
rect 1117 42 1119 48
rect 1156 42 1158 48
rect 1177 42 1179 48
rect 1210 42 1212 48
rect 1231 42 1233 48
rect 1266 42 1268 48
rect 1287 42 1289 48
rect 1320 42 1322 48
rect 1341 42 1343 48
rect 1664 39 1682 41
rect 1655 23 1682 25
rect 1505 -17 1523 -15
rect 1505 -24 1523 -22
rect 1514 -37 1526 -35
rect 1608 -10 1635 -8
rect 1608 -26 1626 -24
rect 1655 -25 1682 -23
rect 1608 -36 1626 -34
rect 1664 -35 1682 -33
rect 1608 -46 1635 -44
rect 1664 -45 1682 -43
rect 1655 -61 1682 -59
rect 1764 -34 1776 -32
rect 1767 -47 1785 -45
rect 1767 -54 1785 -52
rect 132 -116 134 -103
rect 142 -116 144 -103
rect 152 -114 154 -96
rect 219 -116 221 -103
rect 229 -116 231 -103
rect 239 -114 241 -96
rect 312 -116 314 -103
rect 322 -116 324 -103
rect 332 -114 334 -96
rect 552 -112 554 -94
rect 562 -114 564 -101
rect 572 -114 574 -101
rect 645 -112 647 -94
rect 655 -114 657 -101
rect 665 -114 667 -101
rect 732 -112 734 -94
rect 1063 -83 1065 -77
rect 1135 -83 1137 -77
rect 1174 -83 1176 -77
rect 1195 -83 1197 -77
rect 1228 -83 1230 -77
rect 1249 -83 1251 -77
rect 1284 -83 1286 -77
rect 1305 -83 1307 -77
rect 1338 -83 1340 -77
rect 1359 -83 1361 -77
rect 742 -114 744 -101
rect 752 -114 754 -101
rect 1608 -94 1635 -92
rect 1608 -110 1626 -108
rect 1608 -120 1626 -118
rect 1608 -130 1635 -128
rect 54 -170 56 -158
rect 64 -170 66 -160
rect 74 -170 76 -160
rect 140 -169 142 -142
rect 156 -169 158 -151
rect 166 -169 168 -151
rect 176 -169 178 -142
rect 224 -169 226 -142
rect 240 -169 242 -151
rect 250 -169 252 -151
rect 260 -169 262 -142
rect 286 -170 288 -158
rect 296 -170 298 -160
rect 306 -170 308 -160
rect 383 -168 385 -156
rect 393 -168 395 -158
rect 403 -168 405 -158
rect 469 -167 471 -140
rect 485 -167 487 -149
rect 495 -167 497 -149
rect 505 -167 507 -140
rect 553 -167 555 -140
rect 569 -167 571 -149
rect 579 -167 581 -149
rect 589 -167 591 -140
rect 615 -168 617 -156
rect 625 -168 627 -158
rect 635 -168 637 -158
rect 710 -165 712 -153
rect 720 -165 722 -155
rect 730 -165 732 -155
rect 796 -164 798 -137
rect 812 -164 814 -146
rect 822 -164 824 -146
rect 832 -164 834 -137
rect 880 -164 882 -137
rect 896 -164 898 -146
rect 906 -164 908 -146
rect 916 -164 918 -137
rect 1673 -127 1683 -125
rect 1673 -137 1683 -135
rect 942 -165 944 -153
rect 952 -165 954 -155
rect 962 -165 964 -155
rect 1671 -147 1683 -145
rect 1607 -156 1619 -154
rect 1607 -166 1617 -164
rect 1139 -182 1141 -176
rect 1178 -182 1180 -176
rect 1199 -182 1201 -176
rect 1232 -182 1234 -176
rect 1253 -182 1255 -176
rect 1288 -182 1290 -176
rect 1309 -182 1311 -176
rect 1342 -182 1344 -176
rect 1363 -182 1365 -176
rect 1607 -176 1617 -174
rect 147 -272 149 -254
rect 154 -272 156 -254
rect 167 -263 169 -251
rect 1061 -228 1063 -222
rect 1133 -228 1135 -222
rect 1172 -228 1174 -222
rect 1193 -228 1195 -222
rect 1226 -228 1228 -222
rect 1247 -228 1249 -222
rect 1282 -228 1284 -222
rect 1303 -228 1305 -222
rect 1336 -228 1338 -222
rect 1357 -228 1359 -222
rect 476 -270 478 -252
rect 483 -270 485 -252
rect 496 -261 498 -249
rect 803 -267 805 -249
rect 810 -267 812 -249
rect 823 -258 825 -246
rect 1665 -251 1675 -249
rect 1665 -261 1675 -259
rect 53 -316 55 -304
rect 63 -316 65 -306
rect 73 -316 75 -306
rect 139 -315 141 -288
rect 155 -315 157 -297
rect 165 -315 167 -297
rect 175 -315 177 -288
rect 223 -315 225 -288
rect 239 -315 241 -297
rect 249 -315 251 -297
rect 259 -315 261 -288
rect 285 -316 287 -304
rect 295 -316 297 -306
rect 305 -316 307 -306
rect 382 -314 384 -302
rect 392 -314 394 -304
rect 402 -314 404 -304
rect 468 -313 470 -286
rect 484 -313 486 -295
rect 494 -313 496 -295
rect 504 -313 506 -286
rect 552 -313 554 -286
rect 568 -313 570 -295
rect 578 -313 580 -295
rect 588 -313 590 -286
rect 614 -314 616 -302
rect 624 -314 626 -304
rect 634 -314 636 -304
rect 709 -311 711 -299
rect 719 -311 721 -301
rect 729 -311 731 -301
rect 795 -310 797 -283
rect 811 -310 813 -292
rect 821 -310 823 -292
rect 831 -310 833 -283
rect 879 -310 881 -283
rect 895 -310 897 -292
rect 905 -310 907 -292
rect 915 -310 917 -283
rect 941 -311 943 -299
rect 951 -311 953 -301
rect 961 -311 963 -301
rect 1415 -287 1417 -270
rect 1427 -298 1429 -270
rect 1663 -271 1675 -269
rect 1647 -297 1674 -295
rect 1656 -307 1674 -305
rect 1656 -317 1674 -315
rect 1137 -327 1139 -321
rect 1176 -327 1178 -321
rect 1197 -327 1199 -321
rect 1230 -327 1232 -321
rect 1251 -327 1253 -321
rect 1286 -327 1288 -321
rect 1307 -327 1309 -321
rect 1340 -327 1342 -321
rect 1361 -327 1363 -321
rect 146 -418 148 -400
rect 153 -418 155 -400
rect 166 -409 168 -397
rect 1062 -370 1064 -364
rect 1417 -359 1419 -342
rect 1429 -359 1431 -331
rect 1647 -333 1674 -331
rect 1134 -370 1136 -364
rect 1173 -370 1175 -364
rect 1194 -370 1196 -364
rect 1227 -370 1229 -364
rect 1248 -370 1250 -364
rect 1283 -370 1285 -364
rect 1304 -370 1306 -364
rect 1337 -370 1339 -364
rect 1358 -370 1360 -364
rect 475 -416 477 -398
rect 482 -416 484 -398
rect 495 -407 497 -395
rect 802 -413 804 -395
rect 809 -413 811 -395
rect 822 -404 824 -392
rect 1647 -381 1674 -379
rect 1656 -391 1674 -389
rect 1656 -401 1674 -399
rect 1647 -417 1674 -415
rect 347 -463 349 -445
rect 357 -456 359 -443
rect 367 -456 369 -443
rect 440 -463 442 -445
rect 450 -456 452 -443
rect 460 -456 462 -443
rect 527 -463 529 -445
rect 537 -456 539 -443
rect 547 -456 549 -443
rect 1756 -390 1768 -388
rect 1759 -403 1777 -401
rect 1759 -410 1777 -408
rect 1751 -438 1776 -436
rect 1138 -469 1140 -463
rect 1177 -469 1179 -463
rect 1198 -469 1200 -463
rect 1231 -469 1233 -463
rect 1252 -469 1254 -463
rect 1287 -469 1289 -463
rect 1308 -469 1310 -463
rect 1341 -469 1343 -463
rect 1362 -469 1364 -463
rect 1419 -466 1421 -449
rect 1431 -477 1433 -449
rect 1751 -451 1764 -449
rect 1748 -461 1773 -459
rect 1748 -468 1773 -466
rect 1665 -483 1675 -481
rect 1748 -486 1776 -484
rect 1665 -493 1675 -491
rect 1663 -503 1675 -501
rect 1748 -496 1776 -494
rect 1748 -506 1776 -504
<< polycontact >>
rect 1693 465 1697 469
rect 1661 456 1665 460
rect 1685 446 1689 450
rect 1597 433 1601 437
rect 128 415 132 419
rect 138 415 142 419
rect 118 407 122 411
rect 215 415 219 419
rect 225 415 229 419
rect 205 407 209 411
rect 308 415 312 419
rect 318 415 322 419
rect 298 407 302 411
rect 542 417 546 421
rect 552 417 556 421
rect 635 417 639 421
rect 645 417 649 421
rect 562 409 566 413
rect 722 417 726 421
rect 732 417 736 421
rect 655 409 659 413
rect 1040 413 1044 417
rect 1621 423 1625 427
rect 742 409 746 413
rect 1112 412 1116 416
rect 1150 412 1154 416
rect 1171 412 1175 416
rect 1204 412 1208 416
rect 1225 412 1229 416
rect 1260 412 1264 416
rect 1281 412 1285 416
rect 1314 412 1318 416
rect 1335 412 1339 416
rect 1589 414 1593 418
rect 1684 416 1688 420
rect 1684 406 1688 410
rect 1690 385 1694 389
rect 54 352 58 356
rect 115 344 119 348
rect 44 328 48 332
rect 199 344 203 348
rect 152 329 156 333
rect 162 329 166 333
rect 286 352 290 356
rect 383 354 387 358
rect 444 346 448 350
rect 63 320 67 324
rect 131 323 135 327
rect 236 329 240 333
rect 246 329 250 333
rect 276 328 280 332
rect 215 323 219 327
rect 373 330 377 334
rect 295 320 299 324
rect 528 346 532 350
rect 481 331 485 335
rect 491 331 495 335
rect 615 354 619 358
rect 710 357 714 361
rect 771 349 775 353
rect 392 322 396 326
rect 460 325 464 329
rect 565 331 569 335
rect 575 331 579 335
rect 605 330 609 334
rect 544 325 548 329
rect 700 333 704 337
rect 624 322 628 326
rect 855 349 859 353
rect 808 334 812 338
rect 818 334 822 338
rect 942 357 946 361
rect 1669 369 1673 373
rect 1613 362 1617 366
rect 1116 347 1120 351
rect 1154 347 1158 351
rect 1175 347 1179 351
rect 1208 347 1212 351
rect 1229 347 1233 351
rect 1264 347 1268 351
rect 1285 347 1289 351
rect 1318 347 1322 351
rect 1339 347 1343 351
rect 719 325 723 329
rect 787 328 791 332
rect 892 334 896 338
rect 902 334 906 338
rect 932 333 936 337
rect 871 328 875 332
rect 1535 344 1539 348
rect 1527 334 1531 338
rect 1535 332 1539 336
rect 951 325 955 329
rect 1534 324 1538 328
rect 1592 346 1596 350
rect 1598 325 1602 329
rect 1684 332 1688 336
rect 1598 315 1602 319
rect 1684 322 1688 326
rect 133 266 137 270
rect 145 266 149 270
rect 153 265 157 269
rect 462 268 466 272
rect 474 268 478 272
rect 143 258 147 262
rect 482 267 486 271
rect 789 271 793 275
rect 801 271 805 275
rect 472 260 476 264
rect 809 270 813 274
rect 799 263 803 267
rect 1040 268 1044 272
rect 1690 301 1694 305
rect 1748 323 1752 327
rect 1747 315 1751 319
rect 1755 313 1759 317
rect 1747 303 1751 307
rect 1669 285 1673 289
rect 1613 278 1617 282
rect 1112 267 1116 271
rect 1150 267 1154 271
rect 1171 267 1175 271
rect 1204 267 1208 271
rect 1225 267 1229 271
rect 1260 267 1264 271
rect 1281 267 1285 271
rect 1314 267 1318 271
rect 1335 267 1339 271
rect 1380 268 1384 272
rect 1392 268 1396 272
rect 1592 262 1596 266
rect 1598 241 1602 245
rect 53 206 57 210
rect 114 198 118 202
rect 43 182 47 186
rect 198 198 202 202
rect 151 183 155 187
rect 161 183 165 187
rect 285 206 289 210
rect 382 208 386 212
rect 443 200 447 204
rect 62 174 66 178
rect 130 177 134 181
rect 235 183 239 187
rect 245 183 249 187
rect 275 182 279 186
rect 214 177 218 181
rect 372 184 376 188
rect 294 174 298 178
rect 527 200 531 204
rect 480 185 484 189
rect 490 185 494 189
rect 614 208 618 212
rect 709 211 713 215
rect 770 203 774 207
rect 391 176 395 180
rect 459 179 463 183
rect 564 185 568 189
rect 574 185 578 189
rect 604 184 608 188
rect 543 179 547 183
rect 699 187 703 191
rect 623 176 627 180
rect 854 203 858 207
rect 807 188 811 192
rect 817 188 821 192
rect 941 211 945 215
rect 1598 231 1602 235
rect 1693 233 1697 237
rect 1661 224 1665 228
rect 1381 207 1385 211
rect 1393 207 1397 211
rect 1685 214 1689 218
rect 1116 202 1120 206
rect 1154 202 1158 206
rect 1175 202 1179 206
rect 1208 202 1212 206
rect 1229 202 1233 206
rect 1264 202 1268 206
rect 1285 202 1289 206
rect 1318 202 1322 206
rect 1339 202 1343 206
rect 718 179 722 183
rect 786 182 790 186
rect 891 188 895 192
rect 901 188 905 192
rect 931 187 935 191
rect 870 182 874 186
rect 950 179 954 183
rect 1597 201 1601 205
rect 1621 191 1625 195
rect 1589 182 1593 186
rect 132 120 136 124
rect 144 120 148 124
rect 152 119 156 123
rect 461 122 465 126
rect 473 122 477 126
rect 142 112 146 116
rect 481 121 485 125
rect 788 125 792 129
rect 800 125 804 129
rect 471 114 475 118
rect 808 124 812 128
rect 1039 126 1043 130
rect 798 117 802 121
rect 1111 125 1115 129
rect 1149 125 1153 129
rect 1170 125 1174 129
rect 1203 125 1207 129
rect 1224 125 1228 129
rect 1259 125 1263 129
rect 1280 125 1284 129
rect 1313 125 1317 129
rect 1334 125 1338 129
rect 1380 128 1384 132
rect 1392 128 1396 132
rect 1695 105 1699 109
rect 1663 96 1667 100
rect 357 42 361 46
rect 1687 86 1691 90
rect 1599 73 1603 77
rect 337 34 341 38
rect 347 34 351 38
rect 450 42 454 46
rect 1115 60 1119 64
rect 1153 60 1157 64
rect 1174 60 1178 64
rect 1207 60 1211 64
rect 1228 60 1232 64
rect 1263 60 1267 64
rect 1284 60 1288 64
rect 1317 60 1321 64
rect 1338 60 1342 64
rect 430 34 434 38
rect 440 34 444 38
rect 1623 63 1627 67
rect 1591 54 1595 58
rect 1686 56 1690 60
rect 537 42 541 46
rect 1686 46 1690 50
rect 517 34 521 38
rect 527 34 531 38
rect 1692 25 1696 29
rect 1671 9 1675 13
rect 1615 2 1619 6
rect 1537 -16 1541 -12
rect 1529 -26 1533 -22
rect 1537 -28 1541 -24
rect 1536 -36 1540 -32
rect 1594 -14 1598 -10
rect 1600 -35 1604 -31
rect 1686 -28 1690 -24
rect 1600 -45 1604 -41
rect 1686 -38 1690 -34
rect 1692 -59 1696 -55
rect 1750 -37 1754 -33
rect 1749 -45 1753 -41
rect 1757 -47 1761 -43
rect 1749 -57 1753 -53
rect 139 -91 143 -87
rect 149 -91 153 -87
rect 129 -99 133 -95
rect 226 -91 230 -87
rect 236 -91 240 -87
rect 216 -99 220 -95
rect 319 -91 323 -87
rect 329 -91 333 -87
rect 309 -99 313 -95
rect 553 -89 557 -85
rect 563 -89 567 -85
rect 646 -89 650 -85
rect 656 -89 660 -85
rect 573 -97 577 -93
rect 733 -89 737 -85
rect 743 -89 747 -85
rect 666 -97 670 -93
rect 1671 -75 1675 -71
rect 753 -97 757 -93
rect 1061 -98 1065 -94
rect 1615 -82 1619 -78
rect 1133 -99 1137 -95
rect 1171 -99 1175 -95
rect 1192 -99 1196 -95
rect 1225 -99 1229 -95
rect 1246 -99 1250 -95
rect 1281 -99 1285 -95
rect 1302 -99 1306 -95
rect 1335 -99 1339 -95
rect 1356 -99 1360 -95
rect 1594 -98 1598 -94
rect 1600 -119 1604 -115
rect 1600 -129 1604 -125
rect 65 -154 69 -150
rect 126 -162 130 -158
rect 55 -178 59 -174
rect 210 -162 214 -158
rect 163 -177 167 -173
rect 173 -177 177 -173
rect 297 -154 301 -150
rect 394 -152 398 -148
rect 455 -160 459 -156
rect 74 -186 78 -182
rect 142 -183 146 -179
rect 247 -177 251 -173
rect 257 -177 261 -173
rect 287 -178 291 -174
rect 226 -183 230 -179
rect 384 -176 388 -172
rect 306 -186 310 -182
rect 539 -160 543 -156
rect 492 -175 496 -171
rect 502 -175 506 -171
rect 626 -152 630 -148
rect 721 -149 725 -145
rect 782 -157 786 -153
rect 403 -184 407 -180
rect 471 -181 475 -177
rect 576 -175 580 -171
rect 586 -175 590 -171
rect 616 -176 620 -172
rect 555 -181 559 -177
rect 711 -173 715 -169
rect 635 -184 639 -180
rect 866 -157 870 -153
rect 819 -172 823 -168
rect 829 -172 833 -168
rect 1695 -127 1699 -123
rect 1663 -136 1667 -132
rect 953 -149 957 -145
rect 1687 -146 1691 -142
rect 1137 -164 1141 -160
rect 1175 -164 1179 -160
rect 1196 -164 1200 -160
rect 1229 -164 1233 -160
rect 1250 -164 1254 -160
rect 1285 -164 1289 -160
rect 1306 -164 1310 -160
rect 1339 -164 1343 -160
rect 1360 -164 1364 -160
rect 1599 -159 1603 -155
rect 730 -181 734 -177
rect 798 -178 802 -174
rect 903 -172 907 -168
rect 913 -172 917 -168
rect 943 -173 947 -169
rect 882 -178 886 -174
rect 1623 -169 1627 -165
rect 962 -181 966 -177
rect 1591 -178 1595 -174
rect 144 -240 148 -236
rect 156 -240 160 -236
rect 164 -241 168 -237
rect 473 -238 477 -234
rect 485 -238 489 -234
rect 154 -248 158 -244
rect 493 -239 497 -235
rect 800 -235 804 -231
rect 812 -235 816 -231
rect 483 -246 487 -242
rect 820 -236 824 -232
rect 810 -243 814 -239
rect 1059 -243 1063 -239
rect 1131 -244 1135 -240
rect 1169 -244 1173 -240
rect 1190 -244 1194 -240
rect 1223 -244 1227 -240
rect 1244 -244 1248 -240
rect 1279 -244 1283 -240
rect 1300 -244 1304 -240
rect 1333 -244 1337 -240
rect 1354 -244 1358 -240
rect 1687 -251 1691 -247
rect 1412 -266 1416 -262
rect 1424 -266 1428 -262
rect 1655 -260 1659 -256
rect 64 -300 68 -296
rect 125 -308 129 -304
rect 54 -324 58 -320
rect 209 -308 213 -304
rect 162 -323 166 -319
rect 172 -323 176 -319
rect 296 -300 300 -296
rect 393 -298 397 -294
rect 454 -306 458 -302
rect 73 -332 77 -328
rect 141 -329 145 -325
rect 246 -323 250 -319
rect 256 -323 260 -319
rect 286 -324 290 -320
rect 225 -329 229 -325
rect 383 -322 387 -318
rect 305 -332 309 -328
rect 538 -306 542 -302
rect 491 -321 495 -317
rect 501 -321 505 -317
rect 625 -298 629 -294
rect 720 -295 724 -291
rect 781 -303 785 -299
rect 402 -330 406 -326
rect 470 -327 474 -323
rect 575 -321 579 -317
rect 585 -321 589 -317
rect 615 -322 619 -318
rect 554 -327 558 -323
rect 710 -319 714 -315
rect 634 -330 638 -326
rect 865 -303 869 -299
rect 818 -318 822 -314
rect 828 -318 832 -314
rect 952 -295 956 -291
rect 1679 -270 1683 -266
rect 1678 -300 1682 -296
rect 1135 -309 1139 -305
rect 1173 -309 1177 -305
rect 1194 -309 1198 -305
rect 1227 -309 1231 -305
rect 1248 -309 1252 -305
rect 1283 -309 1287 -305
rect 1304 -309 1308 -305
rect 1337 -309 1341 -305
rect 1358 -309 1362 -305
rect 729 -327 733 -323
rect 797 -324 801 -320
rect 902 -318 906 -314
rect 912 -318 916 -314
rect 942 -319 946 -315
rect 881 -324 885 -320
rect 1678 -310 1682 -306
rect 961 -327 965 -323
rect 1684 -331 1688 -327
rect 143 -386 147 -382
rect 155 -386 159 -382
rect 163 -387 167 -383
rect 472 -384 476 -380
rect 484 -384 488 -380
rect 153 -394 157 -390
rect 492 -385 496 -381
rect 1663 -347 1667 -343
rect 1414 -367 1418 -363
rect 1426 -367 1430 -363
rect 799 -381 803 -377
rect 811 -381 815 -377
rect 482 -392 486 -388
rect 819 -382 823 -378
rect 809 -389 813 -385
rect 1060 -385 1064 -381
rect 1132 -386 1136 -382
rect 1170 -386 1174 -382
rect 1191 -386 1195 -382
rect 1224 -386 1228 -382
rect 1245 -386 1249 -382
rect 1280 -386 1284 -382
rect 1301 -386 1305 -382
rect 1334 -386 1338 -382
rect 1355 -386 1359 -382
rect 1678 -384 1682 -380
rect 1678 -394 1682 -390
rect 1684 -415 1688 -411
rect 368 -464 372 -460
rect 348 -472 352 -468
rect 358 -472 362 -468
rect 461 -464 465 -460
rect 1742 -393 1746 -389
rect 1741 -401 1745 -397
rect 1749 -403 1753 -399
rect 1741 -413 1745 -409
rect 1663 -431 1667 -427
rect 1416 -445 1420 -441
rect 1428 -445 1432 -441
rect 1733 -441 1737 -437
rect 1136 -451 1140 -447
rect 1174 -451 1178 -447
rect 1195 -451 1199 -447
rect 1228 -451 1232 -447
rect 1249 -451 1253 -447
rect 1284 -451 1288 -447
rect 1305 -451 1309 -447
rect 1338 -451 1342 -447
rect 1359 -451 1363 -447
rect 1743 -447 1747 -443
rect 441 -472 445 -468
rect 451 -472 455 -468
rect 548 -464 552 -460
rect 528 -472 532 -468
rect 538 -472 542 -468
rect 1740 -461 1744 -457
rect 1687 -483 1691 -479
rect 1740 -480 1744 -476
rect 1655 -492 1659 -488
rect 1740 -487 1744 -483
rect 1679 -502 1683 -498
rect 1740 -497 1744 -493
rect 1740 -507 1744 -503
rect 1769 -572 1773 -568
<< ndcontact >>
rect 1702 468 1706 472
rect 134 441 138 445
rect 221 441 225 445
rect 115 431 119 435
rect 314 441 318 445
rect 145 429 149 433
rect 202 431 206 435
rect 546 443 550 447
rect 232 429 236 433
rect 295 431 299 435
rect 639 443 643 447
rect 325 429 329 433
rect 535 431 539 435
rect 565 433 569 437
rect 726 443 730 447
rect 628 431 632 435
rect 658 433 662 437
rect 715 431 719 435
rect 745 433 749 437
rect 1583 440 1587 444
rect 1711 450 1715 454
rect 1571 429 1575 433
rect 1699 439 1703 443
rect 1027 392 1031 396
rect 1061 392 1065 396
rect 1099 391 1103 395
rect 1580 411 1584 415
rect 1711 423 1715 427
rect 1701 405 1705 409
rect 1133 391 1137 395
rect 1145 392 1149 396
rect 1179 392 1183 396
rect 1199 392 1203 396
rect 1233 392 1237 396
rect 1255 392 1259 396
rect 1289 392 1293 396
rect 1309 392 1313 396
rect 1343 392 1347 396
rect 1699 395 1703 399
rect 1702 383 1706 387
rect 37 314 41 318
rect 115 319 119 323
rect 199 319 203 323
rect 66 311 70 315
rect 129 311 133 315
rect 141 314 145 318
rect 151 312 155 316
rect 48 302 52 306
rect 213 311 217 315
rect 225 314 229 318
rect 235 312 239 316
rect 169 302 173 306
rect 269 314 273 318
rect 366 316 370 320
rect 444 321 448 325
rect 298 311 302 315
rect 528 321 532 325
rect 395 313 399 317
rect 458 313 462 317
rect 470 316 474 320
rect 480 314 484 318
rect 253 302 257 306
rect 280 302 284 306
rect 377 304 381 308
rect 542 313 546 317
rect 554 316 558 320
rect 564 314 568 318
rect 498 304 502 308
rect 598 316 602 320
rect 693 319 697 323
rect 1103 368 1107 372
rect 1137 368 1141 372
rect 1149 367 1153 371
rect 1183 367 1187 371
rect 1203 367 1207 371
rect 1237 367 1241 371
rect 1259 367 1263 371
rect 1293 367 1297 371
rect 1313 367 1317 371
rect 1347 367 1351 371
rect 1694 369 1698 373
rect 1588 362 1592 366
rect 771 324 775 328
rect 627 313 631 317
rect 855 324 859 328
rect 722 316 726 320
rect 785 316 789 320
rect 797 319 801 323
rect 807 317 811 321
rect 582 304 586 308
rect 609 304 613 308
rect 704 307 708 311
rect 869 316 873 320
rect 881 319 885 323
rect 891 317 895 321
rect 825 307 829 311
rect 925 319 929 323
rect 1549 347 1553 351
rect 1549 337 1553 341
rect 1549 327 1553 331
rect 954 316 958 320
rect 1549 317 1553 321
rect 1580 348 1584 352
rect 1583 336 1587 340
rect 1711 339 1715 343
rect 1581 326 1585 330
rect 1701 321 1705 325
rect 909 307 913 311
rect 936 307 940 311
rect 1571 308 1575 312
rect 1699 311 1703 315
rect 130 280 134 284
rect 140 280 144 284
rect 150 280 154 284
rect 160 280 164 284
rect 459 282 463 286
rect 469 282 473 286
rect 479 282 483 286
rect 489 282 493 286
rect 786 285 790 289
rect 796 285 800 289
rect 806 285 810 289
rect 816 285 820 289
rect 1702 299 1706 303
rect 1733 330 1737 334
rect 1733 320 1737 324
rect 1733 310 1737 314
rect 1733 300 1737 304
rect 1694 285 1698 289
rect 1588 278 1592 282
rect 1027 247 1031 251
rect 1061 247 1065 251
rect 1099 246 1103 250
rect 1377 259 1381 263
rect 1133 246 1137 250
rect 1145 247 1149 251
rect 1179 247 1183 251
rect 1199 247 1203 251
rect 1233 247 1237 251
rect 1255 247 1259 251
rect 1289 247 1293 251
rect 1309 247 1313 251
rect 1343 247 1347 251
rect 1388 251 1392 255
rect 1399 259 1403 263
rect 1399 252 1403 256
rect 1580 264 1584 268
rect 1583 252 1587 256
rect 1581 242 1585 246
rect 36 168 40 172
rect 114 173 118 177
rect 198 173 202 177
rect 65 165 69 169
rect 128 165 132 169
rect 140 168 144 172
rect 150 166 154 170
rect 47 156 51 160
rect 212 165 216 169
rect 224 168 228 172
rect 234 166 238 170
rect 168 156 172 160
rect 268 168 272 172
rect 365 170 369 174
rect 443 175 447 179
rect 297 165 301 169
rect 527 175 531 179
rect 394 167 398 171
rect 457 167 461 171
rect 469 170 473 174
rect 479 168 483 172
rect 252 156 256 160
rect 279 156 283 160
rect 376 158 380 162
rect 541 167 545 171
rect 553 170 557 174
rect 563 168 567 172
rect 497 158 501 162
rect 597 170 601 174
rect 692 173 696 177
rect 1103 223 1107 227
rect 1137 223 1141 227
rect 1149 222 1153 226
rect 1183 222 1187 226
rect 1203 222 1207 226
rect 1237 222 1241 226
rect 1259 222 1263 226
rect 1293 222 1297 226
rect 1313 222 1317 226
rect 1347 222 1351 226
rect 1378 216 1382 220
rect 1389 224 1393 228
rect 1400 223 1404 227
rect 1571 224 1575 228
rect 1702 236 1706 240
rect 1400 216 1404 220
rect 1583 208 1587 212
rect 1711 218 1715 222
rect 770 178 774 182
rect 626 167 630 171
rect 854 178 858 182
rect 721 170 725 174
rect 784 170 788 174
rect 796 173 800 177
rect 806 171 810 175
rect 581 158 585 162
rect 608 158 612 162
rect 703 161 707 165
rect 868 170 872 174
rect 880 173 884 177
rect 890 171 894 175
rect 824 161 828 165
rect 924 173 928 177
rect 953 170 957 174
rect 1571 197 1575 201
rect 1699 207 1703 211
rect 1580 179 1584 183
rect 908 161 912 165
rect 935 161 939 165
rect 129 134 133 138
rect 139 134 143 138
rect 149 134 153 138
rect 159 134 163 138
rect 458 136 462 140
rect 468 136 472 140
rect 478 136 482 140
rect 488 136 492 140
rect 785 139 789 143
rect 795 139 799 143
rect 805 139 809 143
rect 815 139 819 143
rect 1026 105 1030 109
rect 1060 105 1064 109
rect 1098 104 1102 108
rect 1377 119 1381 123
rect 1132 104 1136 108
rect 1144 105 1148 109
rect 1178 105 1182 109
rect 1198 105 1202 109
rect 1232 105 1236 109
rect 1254 105 1258 109
rect 1288 105 1292 109
rect 1308 105 1312 109
rect 1388 111 1392 115
rect 1399 119 1403 123
rect 1399 112 1403 116
rect 1342 105 1346 109
rect 1704 108 1708 112
rect 1102 81 1106 85
rect 1136 81 1140 85
rect 1148 80 1152 84
rect 1182 80 1186 84
rect 1202 80 1206 84
rect 1236 80 1240 84
rect 1258 80 1262 84
rect 1292 80 1296 84
rect 1312 80 1316 84
rect 1346 80 1350 84
rect 1585 80 1589 84
rect 1713 90 1717 94
rect 1573 69 1577 73
rect 1701 79 1705 83
rect 1582 51 1586 55
rect 1713 63 1717 67
rect 1703 45 1707 49
rect 1701 35 1705 39
rect 330 20 334 24
rect 360 18 364 22
rect 423 20 427 24
rect 453 18 457 22
rect 510 20 514 24
rect 341 8 345 12
rect 540 18 544 22
rect 434 8 438 12
rect 1704 23 1708 27
rect 521 8 525 12
rect 1696 9 1700 13
rect 1590 2 1594 6
rect 1551 -13 1555 -9
rect 1551 -23 1555 -19
rect 1551 -33 1555 -29
rect 1551 -43 1555 -39
rect 1582 -12 1586 -8
rect 1585 -24 1589 -20
rect 1713 -21 1717 -17
rect 1583 -34 1587 -30
rect 1703 -39 1707 -35
rect 1573 -52 1577 -48
rect 1701 -49 1705 -45
rect 145 -65 149 -61
rect 232 -65 236 -61
rect 126 -75 130 -71
rect 325 -65 329 -61
rect 156 -77 160 -73
rect 213 -75 217 -71
rect 557 -63 561 -59
rect 243 -77 247 -73
rect 306 -75 310 -71
rect 650 -63 654 -59
rect 336 -77 340 -73
rect 546 -75 550 -71
rect 576 -73 580 -69
rect 737 -63 741 -59
rect 639 -75 643 -71
rect 669 -73 673 -69
rect 1704 -61 1708 -57
rect 1735 -30 1739 -26
rect 1735 -40 1739 -36
rect 1735 -50 1739 -46
rect 1735 -60 1739 -56
rect 726 -75 730 -71
rect 756 -73 760 -69
rect 1696 -75 1700 -71
rect 1590 -82 1594 -78
rect 1048 -119 1052 -115
rect 1082 -119 1086 -115
rect 1120 -120 1124 -116
rect 1582 -96 1586 -92
rect 1585 -108 1589 -104
rect 1154 -120 1158 -116
rect 1166 -119 1170 -115
rect 1200 -119 1204 -115
rect 1220 -119 1224 -115
rect 1254 -119 1258 -115
rect 1276 -119 1280 -115
rect 1310 -119 1314 -115
rect 1330 -119 1334 -115
rect 1364 -119 1368 -115
rect 1583 -118 1587 -114
rect 48 -192 52 -188
rect 126 -187 130 -183
rect 210 -187 214 -183
rect 77 -195 81 -191
rect 140 -195 144 -191
rect 152 -192 156 -188
rect 162 -194 166 -190
rect 59 -204 63 -200
rect 224 -195 228 -191
rect 236 -192 240 -188
rect 246 -194 250 -190
rect 180 -204 184 -200
rect 280 -192 284 -188
rect 377 -190 381 -186
rect 455 -185 459 -181
rect 309 -195 313 -191
rect 539 -185 543 -181
rect 406 -193 410 -189
rect 469 -193 473 -189
rect 481 -190 485 -186
rect 491 -192 495 -188
rect 264 -204 268 -200
rect 291 -204 295 -200
rect 388 -202 392 -198
rect 553 -193 557 -189
rect 565 -190 569 -186
rect 575 -192 579 -188
rect 509 -202 513 -198
rect 609 -190 613 -186
rect 704 -187 708 -183
rect 1573 -136 1577 -132
rect 1704 -124 1708 -120
rect 1124 -143 1128 -139
rect 1158 -143 1162 -139
rect 1170 -144 1174 -140
rect 1204 -144 1208 -140
rect 1224 -144 1228 -140
rect 1258 -144 1262 -140
rect 1280 -144 1284 -140
rect 1314 -144 1318 -140
rect 1334 -144 1338 -140
rect 1368 -144 1372 -140
rect 1585 -152 1589 -148
rect 1713 -142 1717 -138
rect 1573 -163 1577 -159
rect 1701 -153 1705 -149
rect 782 -182 786 -178
rect 638 -193 642 -189
rect 866 -182 870 -178
rect 733 -190 737 -186
rect 796 -190 800 -186
rect 808 -187 812 -183
rect 818 -189 822 -185
rect 593 -202 597 -198
rect 620 -202 624 -198
rect 715 -199 719 -195
rect 880 -190 884 -186
rect 892 -187 896 -183
rect 902 -189 906 -185
rect 836 -199 840 -195
rect 936 -187 940 -183
rect 1582 -181 1586 -177
rect 965 -190 969 -186
rect 920 -199 924 -195
rect 947 -199 951 -195
rect 141 -226 145 -222
rect 151 -226 155 -222
rect 161 -226 165 -222
rect 171 -226 175 -222
rect 470 -224 474 -220
rect 480 -224 484 -220
rect 490 -224 494 -220
rect 500 -224 504 -220
rect 797 -221 801 -217
rect 807 -221 811 -217
rect 817 -221 821 -217
rect 827 -221 831 -217
rect 1046 -264 1050 -260
rect 1080 -264 1084 -260
rect 1118 -265 1122 -261
rect 1409 -257 1413 -253
rect 1420 -249 1424 -245
rect 1431 -250 1435 -246
rect 1431 -257 1435 -253
rect 1696 -248 1700 -244
rect 1152 -265 1156 -261
rect 1164 -264 1168 -260
rect 1198 -264 1202 -260
rect 1218 -264 1222 -260
rect 1252 -264 1256 -260
rect 1274 -264 1278 -260
rect 1308 -264 1312 -260
rect 1328 -264 1332 -260
rect 1362 -264 1366 -260
rect 47 -338 51 -334
rect 125 -333 129 -329
rect 209 -333 213 -329
rect 76 -341 80 -337
rect 139 -341 143 -337
rect 151 -338 155 -334
rect 161 -340 165 -336
rect 58 -350 62 -346
rect 223 -341 227 -337
rect 235 -338 239 -334
rect 245 -340 249 -336
rect 179 -350 183 -346
rect 279 -338 283 -334
rect 376 -336 380 -332
rect 454 -331 458 -327
rect 308 -341 312 -337
rect 538 -331 542 -327
rect 405 -339 409 -335
rect 468 -339 472 -335
rect 480 -336 484 -332
rect 490 -338 494 -334
rect 263 -350 267 -346
rect 290 -350 294 -346
rect 387 -348 391 -344
rect 552 -339 556 -335
rect 564 -336 568 -332
rect 574 -338 578 -334
rect 508 -348 512 -344
rect 608 -336 612 -332
rect 703 -333 707 -329
rect 1122 -288 1126 -284
rect 1156 -288 1160 -284
rect 1168 -289 1172 -285
rect 1202 -289 1206 -285
rect 1222 -289 1226 -285
rect 1256 -289 1260 -285
rect 1278 -289 1282 -285
rect 1312 -289 1316 -285
rect 1332 -289 1336 -285
rect 1366 -289 1370 -285
rect 1705 -266 1709 -262
rect 1693 -277 1697 -273
rect 1705 -293 1709 -289
rect 781 -328 785 -324
rect 637 -339 641 -335
rect 865 -328 869 -324
rect 732 -336 736 -332
rect 795 -336 799 -332
rect 807 -333 811 -329
rect 817 -335 821 -331
rect 592 -348 596 -344
rect 619 -348 623 -344
rect 714 -345 718 -341
rect 879 -336 883 -332
rect 891 -333 895 -329
rect 901 -335 905 -331
rect 835 -345 839 -341
rect 935 -333 939 -329
rect 1695 -311 1699 -307
rect 1693 -321 1697 -317
rect 964 -336 968 -332
rect 919 -345 923 -341
rect 946 -345 950 -341
rect 140 -372 144 -368
rect 150 -372 154 -368
rect 160 -372 164 -368
rect 170 -372 174 -368
rect 469 -370 473 -366
rect 479 -370 483 -366
rect 489 -370 493 -366
rect 499 -370 503 -366
rect 796 -367 800 -363
rect 806 -367 810 -363
rect 816 -367 820 -363
rect 826 -367 830 -363
rect 1696 -333 1700 -329
rect 1688 -347 1692 -343
rect 1411 -376 1415 -372
rect 1047 -406 1051 -402
rect 1422 -384 1426 -380
rect 1433 -376 1437 -372
rect 1705 -377 1709 -373
rect 1433 -383 1437 -379
rect 1081 -406 1085 -402
rect 1119 -407 1123 -403
rect 1695 -395 1699 -391
rect 1153 -407 1157 -403
rect 1165 -406 1169 -402
rect 1199 -406 1203 -402
rect 1219 -406 1223 -402
rect 1253 -406 1257 -402
rect 1275 -406 1279 -402
rect 1309 -406 1313 -402
rect 1329 -406 1333 -402
rect 1363 -406 1367 -402
rect 1693 -405 1697 -401
rect 1123 -430 1127 -426
rect 1157 -430 1161 -426
rect 1169 -431 1173 -427
rect 1203 -431 1207 -427
rect 1223 -431 1227 -427
rect 1257 -431 1261 -427
rect 1279 -431 1283 -427
rect 1313 -431 1317 -427
rect 1333 -431 1337 -427
rect 1367 -431 1371 -427
rect 1413 -436 1417 -432
rect 1424 -428 1428 -424
rect 1696 -417 1700 -413
rect 1727 -386 1731 -382
rect 1727 -396 1731 -392
rect 1727 -406 1731 -402
rect 1727 -416 1731 -412
rect 1435 -429 1439 -425
rect 1688 -431 1692 -427
rect 1435 -436 1439 -432
rect 1724 -434 1728 -430
rect 1720 -444 1724 -440
rect 341 -486 345 -482
rect 371 -488 375 -484
rect 434 -486 438 -482
rect 464 -488 468 -484
rect 521 -486 525 -482
rect 352 -498 356 -494
rect 1723 -454 1727 -450
rect 1731 -464 1735 -460
rect 1724 -474 1728 -470
rect 1731 -474 1735 -470
rect 551 -488 555 -484
rect 445 -498 449 -494
rect 1696 -480 1700 -476
rect 1724 -484 1728 -480
rect 532 -498 536 -494
rect 1705 -498 1709 -494
rect 1717 -501 1721 -497
rect 1693 -509 1697 -505
rect 1724 -512 1728 -508
<< pdcontact >>
rect 1672 469 1676 473
rect 1676 459 1680 463
rect 1016 429 1020 433
rect 1060 429 1066 435
rect 1676 449 1680 453
rect 1606 440 1610 444
rect 1676 439 1680 443
rect 1099 429 1103 433
rect 1132 429 1136 433
rect 1145 429 1149 433
rect 1162 429 1166 433
rect 1179 429 1183 433
rect 1199 429 1203 433
rect 1216 429 1220 433
rect 1233 429 1237 433
rect 1255 429 1259 433
rect 1272 429 1276 433
rect 1289 429 1293 433
rect 1309 429 1313 433
rect 1326 429 1330 433
rect 1343 429 1347 433
rect 1606 430 1610 434
rect 115 391 119 395
rect 125 398 129 402
rect 125 391 129 395
rect 135 393 139 397
rect 145 405 149 409
rect 145 398 149 402
rect 202 391 206 395
rect 212 398 216 402
rect 212 391 216 395
rect 222 393 226 397
rect 232 405 236 409
rect 232 398 236 402
rect 295 391 299 395
rect 305 398 309 402
rect 305 391 309 395
rect 315 393 319 397
rect 325 405 329 409
rect 325 398 329 402
rect 535 407 539 411
rect 535 400 539 404
rect 628 407 632 411
rect 545 395 549 399
rect 555 400 559 404
rect 555 393 559 397
rect 628 400 632 404
rect 565 393 569 397
rect 715 407 719 411
rect 638 395 642 399
rect 648 400 652 404
rect 648 393 652 397
rect 715 400 719 404
rect 658 393 662 397
rect 1606 420 1610 424
rect 725 395 729 399
rect 735 400 739 404
rect 735 393 739 397
rect 745 393 749 397
rect 1610 410 1614 414
rect 1660 423 1664 427
rect 1668 413 1672 417
rect 1675 403 1679 407
rect 1654 387 1658 391
rect 1661 387 1665 391
rect 1675 377 1679 381
rect 37 337 41 341
rect 47 337 51 341
rect 57 337 61 341
rect 67 341 71 345
rect 123 338 127 342
rect 133 359 137 363
rect 133 352 137 356
rect 149 338 153 342
rect 159 345 163 349
rect 169 353 173 357
rect 207 338 211 342
rect 217 359 221 363
rect 217 352 221 356
rect 233 338 237 342
rect 243 345 247 349
rect 253 353 257 357
rect 269 337 273 341
rect 279 337 283 341
rect 289 337 293 341
rect 299 341 303 345
rect 366 339 370 343
rect 376 339 380 343
rect 386 339 390 343
rect 396 343 400 347
rect 452 340 456 344
rect 462 361 466 365
rect 462 354 466 358
rect 478 340 482 344
rect 488 347 492 351
rect 498 355 502 359
rect 536 340 540 344
rect 546 361 550 365
rect 546 354 550 358
rect 562 340 566 344
rect 572 347 576 351
rect 582 355 586 359
rect 598 339 602 343
rect 608 339 612 343
rect 618 339 622 343
rect 628 343 632 347
rect 693 342 697 346
rect 703 342 707 346
rect 713 342 717 346
rect 723 346 727 350
rect 779 343 783 347
rect 789 364 793 368
rect 789 357 793 361
rect 805 343 809 347
rect 815 350 819 354
rect 825 358 829 362
rect 863 343 867 347
rect 873 364 877 368
rect 873 357 877 361
rect 889 343 893 347
rect 899 350 903 354
rect 909 358 913 362
rect 925 342 929 346
rect 935 342 939 346
rect 945 342 949 346
rect 955 346 959 350
rect 1511 347 1515 351
rect 1103 330 1107 334
rect 1136 330 1140 334
rect 1149 330 1153 334
rect 1166 330 1170 334
rect 1183 330 1187 334
rect 1203 330 1207 334
rect 1220 330 1224 334
rect 1237 330 1241 334
rect 1259 330 1263 334
rect 1276 330 1280 334
rect 1293 330 1297 334
rect 1313 330 1317 334
rect 1330 330 1334 334
rect 1347 330 1351 334
rect 1504 329 1508 333
rect 1513 317 1517 321
rect 1607 354 1611 358
rect 1621 344 1625 348
rect 1628 344 1632 348
rect 1660 339 1664 343
rect 1607 328 1611 332
rect 1668 329 1672 333
rect 1614 318 1618 322
rect 1675 319 1679 323
rect 1388 302 1392 306
rect 1622 308 1626 312
rect 1016 284 1020 288
rect 130 242 134 246
rect 1060 284 1066 290
rect 1099 284 1103 288
rect 1132 284 1136 288
rect 1145 284 1149 288
rect 1162 284 1166 288
rect 1179 284 1183 288
rect 1199 284 1203 288
rect 1216 284 1220 288
rect 1233 284 1237 288
rect 1255 284 1259 288
rect 1272 284 1276 288
rect 1289 284 1293 288
rect 1309 284 1313 288
rect 1326 284 1330 288
rect 1343 284 1347 288
rect 1377 284 1381 288
rect 1654 303 1658 307
rect 1661 303 1665 307
rect 1399 292 1403 296
rect 1675 293 1679 297
rect 1769 330 1773 334
rect 1778 318 1782 322
rect 1771 300 1775 304
rect 1399 285 1403 289
rect 160 244 164 248
rect 459 244 463 248
rect 148 235 152 239
rect 489 246 493 250
rect 786 247 790 251
rect 477 237 481 241
rect 816 249 820 253
rect 1607 270 1611 274
rect 1621 260 1625 264
rect 1628 260 1632 264
rect 804 240 808 244
rect 1607 244 1611 248
rect 36 191 40 195
rect 46 191 50 195
rect 56 191 60 195
rect 66 195 70 199
rect 122 192 126 196
rect 132 213 136 217
rect 132 206 136 210
rect 148 192 152 196
rect 158 199 162 203
rect 168 207 172 211
rect 206 192 210 196
rect 216 213 220 217
rect 216 206 220 210
rect 232 192 236 196
rect 242 199 246 203
rect 252 207 256 211
rect 268 191 272 195
rect 278 191 282 195
rect 288 191 292 195
rect 298 195 302 199
rect 365 193 369 197
rect 375 193 379 197
rect 385 193 389 197
rect 395 197 399 201
rect 451 194 455 198
rect 461 215 465 219
rect 461 208 465 212
rect 477 194 481 198
rect 487 201 491 205
rect 497 209 501 213
rect 535 194 539 198
rect 545 215 549 219
rect 545 208 549 212
rect 561 194 565 198
rect 571 201 575 205
rect 581 209 585 213
rect 597 193 601 197
rect 607 193 611 197
rect 617 193 621 197
rect 627 197 631 201
rect 692 196 696 200
rect 702 196 706 200
rect 712 196 716 200
rect 722 200 726 204
rect 778 197 782 201
rect 788 218 792 222
rect 788 211 792 215
rect 804 197 808 201
rect 814 204 818 208
rect 824 212 828 216
rect 862 197 866 201
rect 872 218 876 222
rect 872 211 876 215
rect 888 197 892 201
rect 898 204 902 208
rect 908 212 912 216
rect 924 196 928 200
rect 1614 234 1618 238
rect 1622 224 1626 228
rect 1672 237 1676 241
rect 1676 227 1680 231
rect 1676 217 1680 221
rect 1606 208 1610 212
rect 1676 207 1680 211
rect 934 196 938 200
rect 944 196 948 200
rect 954 200 958 204
rect 1378 191 1382 195
rect 1103 185 1107 189
rect 1136 185 1140 189
rect 1149 185 1153 189
rect 1166 185 1170 189
rect 1183 185 1187 189
rect 1203 185 1207 189
rect 1220 185 1224 189
rect 1237 185 1241 189
rect 1259 185 1263 189
rect 1276 185 1280 189
rect 1293 185 1297 189
rect 1313 185 1317 189
rect 1330 185 1334 189
rect 1347 185 1351 189
rect 1389 173 1393 177
rect 1606 198 1610 202
rect 1400 190 1404 194
rect 1606 188 1610 192
rect 1400 183 1404 187
rect 1610 178 1614 182
rect 1388 162 1392 166
rect 1015 142 1019 146
rect 1059 142 1065 148
rect 1098 142 1102 146
rect 1131 142 1135 146
rect 1144 142 1148 146
rect 1161 142 1165 146
rect 1178 142 1182 146
rect 1198 142 1202 146
rect 1215 142 1219 146
rect 1232 142 1236 146
rect 1254 142 1258 146
rect 1271 142 1275 146
rect 1288 142 1292 146
rect 1308 142 1312 146
rect 1325 142 1329 146
rect 1342 142 1346 146
rect 1377 144 1381 148
rect 129 96 133 100
rect 1399 152 1403 156
rect 1399 145 1403 149
rect 159 98 163 102
rect 458 98 462 102
rect 147 89 151 93
rect 488 100 492 104
rect 785 101 789 105
rect 476 91 480 95
rect 815 103 819 107
rect 1674 109 1678 113
rect 803 94 807 98
rect 1678 99 1682 103
rect 330 51 334 55
rect 330 44 334 48
rect 340 56 344 60
rect 350 58 354 62
rect 350 51 354 55
rect 360 58 364 62
rect 423 51 427 55
rect 423 44 427 48
rect 433 56 437 60
rect 443 58 447 62
rect 443 51 447 55
rect 453 58 457 62
rect 1678 89 1682 93
rect 1608 80 1612 84
rect 1678 79 1682 83
rect 1608 70 1612 74
rect 510 51 514 55
rect 510 44 514 48
rect 520 56 524 60
rect 530 58 534 62
rect 530 51 534 55
rect 540 58 544 62
rect 1608 60 1612 64
rect 1612 50 1616 54
rect 1662 63 1666 67
rect 1670 53 1674 57
rect 1102 43 1106 47
rect 1135 43 1139 47
rect 1148 43 1152 47
rect 1165 43 1169 47
rect 1182 43 1186 47
rect 1202 43 1206 47
rect 1219 43 1223 47
rect 1236 43 1240 47
rect 1258 43 1262 47
rect 1275 43 1279 47
rect 1292 43 1296 47
rect 1312 43 1316 47
rect 1329 43 1333 47
rect 1346 43 1350 47
rect 1677 43 1681 47
rect 1656 27 1660 31
rect 1663 27 1667 31
rect 1677 17 1681 21
rect 1513 -13 1517 -9
rect 1506 -31 1510 -27
rect 1515 -43 1519 -39
rect 1609 -6 1613 -2
rect 1623 -16 1627 -12
rect 1630 -16 1634 -12
rect 1662 -21 1666 -17
rect 1609 -32 1613 -28
rect 1670 -31 1674 -27
rect 1616 -42 1620 -38
rect 1677 -41 1681 -37
rect 1624 -52 1628 -48
rect 1656 -57 1660 -53
rect 1663 -57 1667 -53
rect 1677 -67 1681 -63
rect 1771 -30 1775 -26
rect 1780 -42 1784 -38
rect 1773 -60 1777 -56
rect 126 -115 130 -111
rect 136 -108 140 -104
rect 136 -115 140 -111
rect 146 -113 150 -109
rect 156 -101 160 -97
rect 156 -108 160 -104
rect 213 -115 217 -111
rect 223 -108 227 -104
rect 223 -115 227 -111
rect 233 -113 237 -109
rect 243 -101 247 -97
rect 243 -108 247 -104
rect 306 -115 310 -111
rect 316 -108 320 -104
rect 316 -115 320 -111
rect 326 -113 330 -109
rect 336 -101 340 -97
rect 336 -108 340 -104
rect 546 -99 550 -95
rect 546 -106 550 -102
rect 639 -99 643 -95
rect 556 -111 560 -107
rect 566 -106 570 -102
rect 566 -113 570 -109
rect 639 -106 643 -102
rect 576 -113 580 -109
rect 726 -99 730 -95
rect 649 -111 653 -107
rect 659 -106 663 -102
rect 659 -113 663 -109
rect 726 -106 730 -102
rect 669 -113 673 -109
rect 1037 -82 1041 -78
rect 1081 -82 1087 -76
rect 1120 -82 1124 -78
rect 1153 -82 1157 -78
rect 1166 -82 1170 -78
rect 1183 -82 1187 -78
rect 1200 -82 1204 -78
rect 1220 -82 1224 -78
rect 1237 -82 1241 -78
rect 1254 -82 1258 -78
rect 1276 -82 1280 -78
rect 1293 -82 1297 -78
rect 1310 -82 1314 -78
rect 1330 -82 1334 -78
rect 1347 -82 1351 -78
rect 1364 -82 1368 -78
rect 736 -111 740 -107
rect 746 -106 750 -102
rect 746 -113 750 -109
rect 756 -113 760 -109
rect 1609 -90 1613 -86
rect 1623 -100 1627 -96
rect 1630 -100 1634 -96
rect 1609 -116 1613 -112
rect 1616 -126 1620 -122
rect 48 -169 52 -165
rect 58 -169 62 -165
rect 68 -169 72 -165
rect 78 -165 82 -161
rect 134 -168 138 -164
rect 144 -147 148 -143
rect 144 -154 148 -150
rect 160 -168 164 -164
rect 170 -161 174 -157
rect 180 -153 184 -149
rect 218 -168 222 -164
rect 228 -147 232 -143
rect 228 -154 232 -150
rect 244 -168 248 -164
rect 254 -161 258 -157
rect 264 -153 268 -149
rect 280 -169 284 -165
rect 290 -169 294 -165
rect 300 -169 304 -165
rect 310 -165 314 -161
rect 377 -167 381 -163
rect 387 -167 391 -163
rect 397 -167 401 -163
rect 407 -163 411 -159
rect 463 -166 467 -162
rect 473 -145 477 -141
rect 473 -152 477 -148
rect 489 -166 493 -162
rect 499 -159 503 -155
rect 509 -151 513 -147
rect 547 -166 551 -162
rect 557 -145 561 -141
rect 557 -152 561 -148
rect 573 -166 577 -162
rect 583 -159 587 -155
rect 593 -151 597 -147
rect 609 -167 613 -163
rect 619 -167 623 -163
rect 629 -167 633 -163
rect 639 -163 643 -159
rect 704 -164 708 -160
rect 714 -164 718 -160
rect 724 -164 728 -160
rect 734 -160 738 -156
rect 790 -163 794 -159
rect 800 -142 804 -138
rect 800 -149 804 -145
rect 816 -163 820 -159
rect 826 -156 830 -152
rect 836 -148 840 -144
rect 874 -163 878 -159
rect 884 -142 888 -138
rect 884 -149 888 -145
rect 900 -163 904 -159
rect 910 -156 914 -152
rect 1624 -136 1628 -132
rect 1674 -123 1678 -119
rect 1678 -133 1682 -129
rect 920 -148 924 -144
rect 936 -164 940 -160
rect 946 -164 950 -160
rect 956 -164 960 -160
rect 966 -160 970 -156
rect 1678 -143 1682 -139
rect 1608 -152 1612 -148
rect 1678 -153 1682 -149
rect 1608 -162 1612 -158
rect 1608 -172 1612 -168
rect 1124 -181 1128 -177
rect 1157 -181 1161 -177
rect 1170 -181 1174 -177
rect 1187 -181 1191 -177
rect 1204 -181 1208 -177
rect 1224 -181 1228 -177
rect 1241 -181 1245 -177
rect 1258 -181 1262 -177
rect 1280 -181 1284 -177
rect 1297 -181 1301 -177
rect 1314 -181 1318 -177
rect 1334 -181 1338 -177
rect 1351 -181 1355 -177
rect 1368 -181 1372 -177
rect 1612 -182 1616 -178
rect 141 -264 145 -260
rect 1035 -227 1039 -223
rect 1079 -227 1085 -221
rect 1118 -227 1122 -223
rect 1151 -227 1155 -223
rect 1164 -227 1168 -223
rect 1181 -227 1185 -223
rect 1198 -227 1202 -223
rect 1218 -227 1222 -223
rect 1235 -227 1239 -223
rect 1252 -227 1256 -223
rect 1274 -227 1278 -223
rect 1291 -227 1295 -223
rect 1308 -227 1312 -223
rect 1328 -227 1332 -223
rect 1345 -227 1349 -223
rect 1362 -227 1366 -223
rect 171 -262 175 -258
rect 470 -262 474 -258
rect 159 -271 163 -267
rect 500 -260 504 -256
rect 797 -259 801 -255
rect 488 -269 492 -265
rect 827 -257 831 -253
rect 815 -266 819 -262
rect 1666 -247 1670 -243
rect 1670 -257 1674 -253
rect 47 -315 51 -311
rect 57 -315 61 -311
rect 67 -315 71 -311
rect 77 -311 81 -307
rect 133 -314 137 -310
rect 143 -293 147 -289
rect 143 -300 147 -296
rect 159 -314 163 -310
rect 169 -307 173 -303
rect 179 -299 183 -295
rect 217 -314 221 -310
rect 227 -293 231 -289
rect 227 -300 231 -296
rect 243 -314 247 -310
rect 253 -307 257 -303
rect 263 -299 267 -295
rect 279 -315 283 -311
rect 289 -315 293 -311
rect 299 -315 303 -311
rect 309 -311 313 -307
rect 376 -313 380 -309
rect 386 -313 390 -309
rect 396 -313 400 -309
rect 406 -309 410 -305
rect 462 -312 466 -308
rect 472 -291 476 -287
rect 472 -298 476 -294
rect 488 -312 492 -308
rect 498 -305 502 -301
rect 508 -297 512 -293
rect 546 -312 550 -308
rect 556 -291 560 -287
rect 556 -298 560 -294
rect 572 -312 576 -308
rect 582 -305 586 -301
rect 592 -297 596 -293
rect 608 -313 612 -309
rect 618 -313 622 -309
rect 628 -313 632 -309
rect 638 -309 642 -305
rect 703 -310 707 -306
rect 713 -310 717 -306
rect 723 -310 727 -306
rect 733 -306 737 -302
rect 789 -309 793 -305
rect 799 -288 803 -284
rect 799 -295 803 -291
rect 815 -309 819 -305
rect 825 -302 829 -298
rect 835 -294 839 -290
rect 873 -309 877 -305
rect 883 -288 887 -284
rect 883 -295 887 -291
rect 899 -309 903 -305
rect 909 -302 913 -298
rect 1409 -282 1413 -278
rect 919 -294 923 -290
rect 935 -310 939 -306
rect 945 -310 949 -306
rect 955 -310 959 -306
rect 965 -306 969 -302
rect 1420 -300 1424 -296
rect 1670 -267 1674 -263
rect 1670 -277 1674 -273
rect 1431 -283 1435 -279
rect 1431 -290 1435 -286
rect 1654 -293 1658 -289
rect 1662 -303 1666 -299
rect 1669 -313 1673 -309
rect 1122 -326 1126 -322
rect 1155 -326 1159 -322
rect 1168 -326 1172 -322
rect 1185 -326 1189 -322
rect 1202 -326 1206 -322
rect 1222 -326 1226 -322
rect 1239 -326 1243 -322
rect 1256 -326 1260 -322
rect 1278 -326 1282 -322
rect 1295 -326 1299 -322
rect 1312 -326 1316 -322
rect 1332 -326 1336 -322
rect 1349 -326 1353 -322
rect 1366 -326 1370 -322
rect 1422 -333 1426 -329
rect 1648 -329 1652 -325
rect 1655 -329 1659 -325
rect 1411 -351 1415 -347
rect 140 -410 144 -406
rect 1036 -369 1040 -365
rect 1080 -369 1086 -363
rect 1433 -343 1437 -339
rect 1669 -339 1673 -335
rect 1433 -350 1437 -346
rect 1119 -369 1123 -365
rect 1152 -369 1156 -365
rect 1165 -369 1169 -365
rect 1182 -369 1186 -365
rect 1199 -369 1203 -365
rect 1219 -369 1223 -365
rect 1236 -369 1240 -365
rect 1253 -369 1257 -365
rect 1275 -369 1279 -365
rect 1292 -369 1296 -365
rect 1309 -369 1313 -365
rect 1329 -369 1333 -365
rect 1346 -369 1350 -365
rect 1363 -369 1367 -365
rect 170 -408 174 -404
rect 469 -408 473 -404
rect 158 -417 162 -413
rect 499 -406 503 -402
rect 796 -405 800 -401
rect 487 -415 491 -411
rect 826 -403 830 -399
rect 1654 -377 1658 -373
rect 814 -412 818 -408
rect 1662 -387 1666 -383
rect 1669 -397 1673 -393
rect 1648 -413 1652 -409
rect 1655 -413 1659 -409
rect 341 -455 345 -451
rect 341 -462 345 -458
rect 351 -450 355 -446
rect 361 -448 365 -444
rect 361 -455 365 -451
rect 371 -448 375 -444
rect 434 -455 438 -451
rect 434 -462 438 -458
rect 444 -450 448 -446
rect 454 -448 458 -444
rect 454 -455 458 -451
rect 464 -448 468 -444
rect 521 -455 525 -451
rect 521 -462 525 -458
rect 531 -450 535 -446
rect 541 -448 545 -444
rect 541 -455 545 -451
rect 551 -448 555 -444
rect 1669 -423 1673 -419
rect 1763 -386 1767 -382
rect 1772 -398 1776 -394
rect 1765 -416 1769 -412
rect 1752 -434 1756 -430
rect 1759 -434 1763 -430
rect 1413 -461 1417 -457
rect 1123 -468 1127 -464
rect 1156 -468 1160 -464
rect 1169 -468 1173 -464
rect 1186 -468 1190 -464
rect 1203 -468 1207 -464
rect 1223 -468 1227 -464
rect 1240 -468 1244 -464
rect 1257 -468 1261 -464
rect 1279 -468 1283 -464
rect 1296 -468 1300 -464
rect 1313 -468 1317 -464
rect 1333 -468 1337 -464
rect 1350 -468 1354 -464
rect 1367 -468 1371 -464
rect 1424 -479 1428 -475
rect 1772 -445 1776 -441
rect 1435 -462 1439 -458
rect 1435 -469 1439 -465
rect 1752 -457 1756 -453
rect 1666 -479 1670 -475
rect 1670 -489 1674 -485
rect 1764 -480 1768 -476
rect 1771 -480 1775 -476
rect 1756 -492 1760 -488
rect 1763 -492 1767 -488
rect 1670 -499 1674 -495
rect 1764 -502 1768 -498
rect 1771 -502 1775 -498
rect 1670 -509 1674 -505
rect 1749 -512 1753 -508
rect 1756 -512 1760 -508
<< m2contact >>
rect 474 457 479 463
rect 110 448 115 453
rect 463 451 467 455
rect 946 450 951 455
rect 999 441 1003 445
rect 462 436 467 441
rect 498 436 503 441
rect 32 430 37 436
rect 110 424 114 428
rect 102 398 107 403
rect 198 424 202 428
rect 194 398 198 402
rect 291 424 295 428
rect 339 429 343 433
rect 515 429 520 434
rect 243 397 247 401
rect 287 398 291 402
rect 980 437 984 441
rect 412 417 417 422
rect 473 418 478 423
rect 569 426 573 430
rect 339 406 343 410
rect 516 406 521 411
rect 573 400 577 404
rect 339 389 343 393
rect 517 389 521 393
rect 604 399 608 404
rect 662 425 666 429
rect 1025 441 1029 445
rect 749 425 753 429
rect 666 400 670 404
rect 679 402 683 406
rect 232 372 236 376
rect 269 373 274 377
rect 580 378 585 383
rect 615 378 619 383
rect 678 378 682 382
rect 692 377 696 381
rect 702 402 706 406
rect 944 408 950 414
rect 1047 414 1051 418
rect 1119 413 1123 417
rect 754 400 759 404
rect 702 378 706 382
rect 1062 404 1066 408
rect 1122 403 1126 407
rect 1144 413 1148 417
rect 1166 414 1170 418
rect 1134 403 1138 407
rect 1186 421 1190 425
rect 1196 413 1200 417
rect 1163 399 1167 403
rect 1220 404 1224 408
rect 1253 413 1257 417
rect 1289 416 1293 420
rect 1252 405 1256 409
rect 1269 408 1273 412
rect 1279 406 1283 410
rect 1242 398 1246 402
rect 1328 414 1332 418
rect 1342 407 1346 411
rect 1311 399 1315 403
rect 60 352 64 356
rect 203 352 207 356
rect 36 324 40 328
rect 68 326 72 330
rect 105 326 109 330
rect 125 325 129 329
rect 261 343 265 347
rect 172 325 176 329
rect 209 325 213 329
rect 292 352 296 356
rect 307 343 311 347
rect 322 343 326 347
rect 261 309 265 313
rect 300 327 304 331
rect 17 298 21 302
rect 302 299 308 305
rect 129 257 133 261
rect 120 249 124 253
rect 322 275 326 279
rect 389 354 393 358
rect 418 345 422 350
rect 365 326 369 330
rect 397 328 401 332
rect 410 314 414 319
rect 532 354 536 358
rect 434 328 438 332
rect 454 327 458 331
rect 589 347 593 351
rect 501 327 505 331
rect 538 327 542 331
rect 621 354 625 358
rect 590 311 594 315
rect 629 329 633 333
rect 342 298 349 305
rect 629 301 635 307
rect 579 287 584 292
rect 347 275 351 279
rect 419 275 423 279
rect 458 259 462 263
rect 449 251 453 255
rect 641 272 645 276
rect 302 227 307 231
rect 322 226 327 231
rect 59 206 63 210
rect 716 357 720 361
rect 859 357 863 361
rect 751 347 755 351
rect 692 329 696 333
rect 724 331 728 335
rect 761 331 765 335
rect 781 330 785 334
rect 836 349 840 353
rect 828 330 832 334
rect 752 314 756 318
rect 837 314 841 318
rect 914 350 919 354
rect 865 330 869 334
rect 948 357 952 361
rect 917 314 921 318
rect 956 332 960 336
rect 1138 356 1142 360
rect 1086 350 1091 355
rect 669 300 676 307
rect 753 284 758 289
rect 673 272 677 276
rect 744 272 748 276
rect 766 277 770 281
rect 785 262 789 266
rect 776 254 780 258
rect 829 277 833 281
rect 837 271 841 276
rect 766 246 770 250
rect 754 240 758 244
rect 836 236 841 243
rect 1123 346 1127 350
rect 1224 355 1228 359
rect 1256 354 1260 358
rect 1148 346 1152 350
rect 1170 346 1174 350
rect 1200 346 1204 350
rect 1283 353 1287 357
rect 1257 346 1261 350
rect 1315 360 1319 364
rect 1346 352 1350 356
rect 1293 343 1297 347
rect 1332 345 1336 349
rect 1190 338 1194 342
rect 1084 317 1089 322
rect 1686 470 1690 474
rect 1559 463 1563 467
rect 1661 462 1665 466
rect 1593 441 1597 445
rect 1560 367 1564 371
rect 1621 417 1625 421
rect 1676 429 1680 433
rect 1704 431 1708 435
rect 1595 409 1599 413
rect 1580 395 1585 400
rect 1621 395 1625 399
rect 1595 372 1599 376
rect 1518 357 1522 361
rect 1526 348 1530 352
rect 1594 352 1598 356
rect 1688 379 1692 383
rect 1661 373 1665 377
rect 1660 353 1664 357
rect 1703 354 1707 358
rect 1108 299 1112 303
rect 1047 269 1051 273
rect 1119 268 1123 272
rect 1062 259 1066 263
rect 1144 268 1148 272
rect 1166 268 1170 272
rect 1186 276 1190 280
rect 1196 268 1200 272
rect 1134 258 1138 262
rect 1220 259 1224 263
rect 1253 268 1257 272
rect 1289 271 1293 275
rect 1252 260 1256 264
rect 1269 263 1273 267
rect 1279 261 1283 265
rect 1242 253 1246 257
rect 1328 269 1332 273
rect 1342 262 1346 266
rect 1311 254 1315 258
rect 955 236 959 240
rect 35 178 39 182
rect 67 180 71 184
rect 104 180 108 184
rect 124 179 128 183
rect 171 179 175 183
rect 202 206 206 210
rect 291 206 295 210
rect 308 198 312 202
rect 208 179 212 183
rect 260 187 264 191
rect 185 163 189 167
rect 260 163 264 167
rect 299 181 303 185
rect 302 153 310 160
rect 251 143 255 147
rect 321 144 325 148
rect 128 111 132 115
rect 119 103 123 107
rect 246 124 252 130
rect 275 124 280 129
rect 300 124 305 129
rect 321 124 326 129
rect 388 208 392 212
rect 531 208 535 212
rect 424 189 428 193
rect 364 180 368 184
rect 396 182 400 186
rect 433 182 437 186
rect 453 181 457 185
rect 500 181 504 185
rect 424 165 428 169
rect 589 193 593 197
rect 620 208 624 212
rect 537 181 541 185
rect 589 165 593 169
rect 628 183 632 187
rect 339 153 344 158
rect 629 154 633 158
rect 348 144 352 148
rect 424 139 428 143
rect 424 121 428 125
rect 383 91 387 95
rect 457 113 461 117
rect 448 105 452 109
rect 514 131 520 136
rect 602 131 607 136
rect 497 98 502 103
rect 396 91 400 95
rect 385 77 389 81
rect 407 77 411 81
rect 585 76 589 81
rect 396 62 400 66
rect 368 25 373 30
rect 388 14 392 18
rect 498 54 502 59
rect 465 42 469 47
rect 461 25 466 30
rect 554 42 558 46
rect 715 211 719 215
rect 858 211 862 215
rect 691 183 695 187
rect 723 185 727 189
rect 760 185 764 189
rect 780 184 784 188
rect 827 184 831 188
rect 916 195 920 199
rect 947 211 951 215
rect 864 184 868 188
rect 916 168 920 172
rect 955 186 959 190
rect 669 154 673 158
rect 727 145 731 149
rect 666 131 671 136
rect 700 131 705 136
rect 784 116 788 120
rect 775 108 779 112
rect 832 133 838 138
rect 727 104 731 108
rect 1348 238 1352 242
rect 1138 211 1142 215
rect 1123 201 1127 205
rect 1224 210 1228 214
rect 1256 209 1260 213
rect 1148 201 1152 205
rect 1170 201 1174 205
rect 1200 201 1204 205
rect 1283 208 1287 212
rect 1257 201 1261 205
rect 1315 215 1319 219
rect 1346 207 1350 211
rect 1293 198 1297 202
rect 1332 200 1336 204
rect 1190 193 1194 197
rect 1419 302 1426 308
rect 1370 277 1374 281
rect 1519 307 1523 311
rect 1514 290 1521 296
rect 1594 305 1598 309
rect 1688 342 1692 346
rect 1725 353 1729 357
rect 1369 239 1373 243
rect 1426 235 1431 241
rect 1372 198 1376 202
rect 1404 199 1408 203
rect 1050 158 1054 162
rect 1105 154 1109 158
rect 1046 127 1050 131
rect 1118 126 1122 130
rect 1061 117 1065 121
rect 1143 126 1147 130
rect 1165 126 1169 130
rect 1185 134 1189 138
rect 1195 126 1199 130
rect 1133 116 1137 120
rect 1219 117 1223 121
rect 1252 126 1256 130
rect 1288 129 1292 133
rect 1251 118 1255 122
rect 1268 121 1272 125
rect 1278 119 1282 123
rect 1241 111 1245 115
rect 1327 127 1331 131
rect 1341 120 1345 124
rect 1310 112 1314 116
rect 677 69 682 75
rect 1007 48 1011 52
rect 1009 38 1015 44
rect 990 34 994 38
rect 546 25 551 30
rect 999 26 1003 30
rect 1137 69 1141 73
rect 1122 59 1126 63
rect 1059 45 1063 49
rect 1223 68 1227 72
rect 1255 67 1259 71
rect 1147 59 1151 63
rect 1169 59 1173 63
rect 1199 59 1203 63
rect 1282 66 1286 70
rect 1256 59 1260 63
rect 1314 73 1318 77
rect 1345 65 1349 69
rect 1292 56 1296 60
rect 1331 58 1335 62
rect 1189 51 1193 55
rect 1058 30 1062 34
rect 1091 29 1096 33
rect 1353 29 1357 33
rect 1372 127 1376 131
rect 1403 132 1407 136
rect 1395 91 1400 95
rect 1621 274 1625 278
rect 1594 268 1598 272
rect 1551 239 1556 244
rect 1540 229 1545 234
rect 1510 203 1515 208
rect 1511 189 1516 194
rect 1559 226 1563 230
rect 1559 204 1563 208
rect 1688 295 1692 299
rect 1756 299 1760 303
rect 1764 290 1768 294
rect 1687 275 1691 279
rect 1687 238 1691 242
rect 1578 216 1582 220
rect 1604 216 1608 220
rect 1661 230 1665 234
rect 1744 254 1748 258
rect 1772 252 1777 256
rect 1689 206 1693 210
rect 1621 185 1625 189
rect 1717 183 1725 191
rect 1596 177 1600 181
rect 1510 143 1515 148
rect 1725 157 1729 161
rect 1690 138 1697 144
rect 1521 127 1526 132
rect 1547 128 1552 133
rect 1379 19 1384 23
rect 182 0 187 7
rect 312 3 319 10
rect 1048 5 1053 10
rect 1415 19 1419 23
rect 976 -26 983 -21
rect 998 -26 1004 -20
rect 485 -49 490 -43
rect 121 -58 126 -53
rect 43 -76 48 -70
rect 121 -82 125 -78
rect 113 -108 118 -103
rect 209 -82 213 -78
rect 205 -108 209 -104
rect 302 -82 306 -78
rect 350 -77 354 -73
rect 423 -77 429 -71
rect 526 -77 531 -72
rect 254 -109 258 -105
rect 298 -108 302 -104
rect 431 -87 435 -82
rect 484 -88 489 -83
rect 350 -100 354 -96
rect 411 -99 417 -93
rect 580 -80 584 -76
rect 527 -99 532 -95
rect 392 -110 398 -104
rect 486 -109 491 -104
rect 513 -109 518 -104
rect 584 -106 588 -102
rect 350 -117 354 -113
rect 528 -117 532 -113
rect 615 -107 619 -102
rect 673 -81 677 -77
rect 760 -81 764 -77
rect 1019 -11 1023 -7
rect 1053 -18 1057 -14
rect 1109 -16 1114 -11
rect 1014 -26 1021 -18
rect 1131 -27 1139 -20
rect 1099 -38 1104 -34
rect 1107 -72 1112 -67
rect 677 -106 681 -102
rect 690 -104 694 -100
rect 243 -134 247 -130
rect 280 -133 285 -129
rect 591 -128 596 -123
rect 626 -128 630 -123
rect 689 -128 693 -124
rect 703 -129 707 -125
rect 713 -104 717 -100
rect 990 -95 994 -90
rect 1039 -95 1044 -91
rect 1068 -97 1072 -93
rect 765 -106 770 -102
rect 1140 -98 1144 -94
rect 1083 -107 1087 -103
rect 1165 -98 1169 -94
rect 1187 -98 1191 -94
rect 1207 -90 1211 -86
rect 1217 -98 1221 -94
rect 1155 -108 1159 -104
rect 1241 -107 1245 -103
rect 1274 -98 1278 -94
rect 1310 -95 1314 -91
rect 1273 -106 1277 -102
rect 1290 -103 1294 -99
rect 1300 -105 1304 -101
rect 1263 -113 1267 -109
rect 1349 -97 1353 -93
rect 1363 -104 1367 -100
rect 1332 -112 1336 -108
rect 713 -128 717 -124
rect 71 -154 75 -150
rect 214 -154 218 -150
rect 47 -182 51 -178
rect 79 -180 83 -176
rect 116 -180 120 -176
rect 136 -181 140 -177
rect 183 -181 187 -177
rect 303 -153 307 -149
rect 317 -162 321 -158
rect 220 -181 224 -177
rect 272 -173 276 -169
rect 272 -197 276 -193
rect 311 -179 315 -175
rect 28 -208 32 -204
rect 313 -207 319 -201
rect 302 -221 307 -216
rect 140 -249 144 -245
rect 131 -257 135 -253
rect 333 -231 337 -227
rect 400 -152 404 -148
rect 543 -152 547 -148
rect 376 -180 380 -176
rect 408 -178 412 -174
rect 445 -178 449 -174
rect 465 -179 469 -175
rect 600 -159 604 -155
rect 512 -179 516 -175
rect 549 -179 553 -175
rect 632 -152 636 -148
rect 601 -195 605 -191
rect 640 -177 644 -173
rect 353 -208 360 -201
rect 640 -205 646 -199
rect 444 -219 449 -214
rect 358 -231 362 -227
rect 430 -231 434 -227
rect 301 -259 306 -253
rect 333 -259 337 -254
rect 540 -219 545 -214
rect 629 -219 634 -215
rect 469 -247 473 -243
rect 443 -259 448 -254
rect 460 -255 464 -251
rect 652 -234 656 -230
rect 629 -251 633 -247
rect 727 -149 731 -145
rect 870 -149 874 -145
rect 762 -159 766 -155
rect 747 -167 751 -163
rect 703 -177 707 -173
rect 735 -175 739 -171
rect 745 -191 749 -186
rect 772 -175 776 -171
rect 792 -176 796 -172
rect 847 -157 851 -153
rect 839 -176 843 -172
rect 763 -192 767 -188
rect 848 -192 852 -188
rect 925 -156 930 -152
rect 876 -176 880 -172
rect 959 -149 963 -145
rect 928 -192 932 -188
rect 967 -174 971 -170
rect 680 -206 687 -199
rect 313 -279 318 -275
rect 333 -280 338 -275
rect 70 -300 74 -296
rect 46 -328 50 -324
rect 78 -326 82 -322
rect 115 -326 119 -322
rect 135 -327 139 -323
rect 182 -327 186 -323
rect 213 -300 217 -296
rect 271 -312 275 -308
rect 219 -327 223 -323
rect 196 -343 200 -339
rect 302 -300 306 -296
rect 318 -308 322 -304
rect 333 -308 337 -304
rect 271 -343 275 -339
rect 310 -325 314 -321
rect 313 -353 321 -346
rect 262 -363 266 -359
rect 139 -395 143 -391
rect 130 -403 134 -399
rect 257 -382 263 -376
rect 286 -382 291 -377
rect 293 -406 297 -402
rect 311 -382 316 -377
rect 332 -382 337 -377
rect 399 -298 403 -294
rect 542 -298 546 -294
rect 435 -317 439 -313
rect 375 -326 379 -322
rect 407 -324 411 -320
rect 444 -324 448 -320
rect 464 -325 468 -321
rect 511 -325 515 -321
rect 435 -341 439 -337
rect 600 -314 604 -310
rect 631 -298 635 -294
rect 548 -325 552 -321
rect 600 -341 604 -337
rect 639 -323 643 -319
rect 350 -353 355 -348
rect 640 -352 644 -348
rect 384 -361 388 -356
rect 446 -359 450 -355
rect 435 -367 439 -363
rect 359 -374 363 -369
rect 411 -374 415 -369
rect 384 -383 389 -377
rect 588 -359 592 -355
rect 312 -406 317 -401
rect 332 -406 337 -401
rect 385 -416 389 -411
rect 435 -385 439 -381
rect 468 -393 472 -389
rect 459 -401 463 -397
rect 525 -375 531 -370
rect 613 -375 618 -370
rect 632 -394 637 -390
rect 508 -408 513 -403
rect 407 -415 411 -411
rect 712 -225 717 -220
rect 764 -222 769 -217
rect 684 -234 688 -230
rect 755 -234 759 -230
rect 777 -229 781 -225
rect 796 -244 800 -240
rect 787 -252 791 -248
rect 840 -229 844 -225
rect 848 -235 852 -230
rect 777 -260 781 -256
rect 696 -267 700 -262
rect 765 -266 769 -262
rect 847 -270 852 -263
rect 960 -272 964 -267
rect 1019 -147 1025 -141
rect 1159 -155 1163 -151
rect 1144 -165 1148 -161
rect 1245 -156 1249 -152
rect 1277 -157 1281 -153
rect 1169 -165 1173 -161
rect 1191 -165 1195 -161
rect 1221 -165 1225 -161
rect 1304 -158 1308 -154
rect 1278 -165 1282 -161
rect 1336 -151 1340 -147
rect 1367 -159 1371 -155
rect 1314 -168 1318 -164
rect 1353 -166 1357 -162
rect 1211 -173 1215 -169
rect 1019 -192 1025 -186
rect 1406 -147 1412 -141
rect 1128 -212 1132 -208
rect 1066 -242 1070 -238
rect 1138 -243 1142 -239
rect 1081 -252 1085 -248
rect 1163 -243 1167 -239
rect 1185 -243 1189 -239
rect 1205 -235 1209 -231
rect 1215 -243 1219 -239
rect 1153 -253 1157 -249
rect 1239 -252 1243 -248
rect 1272 -243 1276 -239
rect 1308 -240 1312 -236
rect 1271 -251 1275 -247
rect 1288 -248 1292 -244
rect 1298 -250 1302 -246
rect 1261 -258 1265 -254
rect 1347 -242 1351 -238
rect 1361 -249 1365 -245
rect 1330 -257 1334 -253
rect 726 -295 730 -291
rect 751 -304 755 -299
rect 702 -323 706 -319
rect 734 -321 738 -317
rect 869 -295 873 -291
rect 771 -321 775 -317
rect 791 -322 795 -318
rect 838 -322 842 -318
rect 749 -334 753 -329
rect 927 -311 931 -307
rect 958 -295 962 -291
rect 875 -322 879 -318
rect 927 -338 931 -334
rect 966 -320 970 -316
rect 680 -352 684 -348
rect 738 -361 742 -357
rect 677 -375 682 -370
rect 711 -375 716 -370
rect 738 -402 742 -398
rect 754 -383 758 -379
rect 843 -373 849 -368
rect 795 -390 799 -386
rect 786 -398 790 -394
rect 753 -407 757 -402
rect 1368 -279 1372 -275
rect 1322 -286 1326 -282
rect 1157 -300 1161 -296
rect 1142 -310 1146 -306
rect 1243 -301 1247 -297
rect 1275 -302 1279 -298
rect 1167 -310 1171 -306
rect 1189 -310 1193 -306
rect 1219 -310 1223 -306
rect 1302 -303 1306 -299
rect 1276 -310 1280 -306
rect 1312 -313 1316 -309
rect 1209 -318 1213 -314
rect 1334 -296 1338 -292
rect 1365 -304 1369 -300
rect 1351 -311 1355 -307
rect 1521 98 1525 102
rect 1537 101 1541 105
rect 1537 75 1541 79
rect 1688 110 1692 114
rect 1663 102 1667 106
rect 1724 117 1729 121
rect 1595 81 1599 85
rect 1552 60 1556 64
rect 1623 57 1627 61
rect 1678 71 1682 75
rect 1706 71 1710 75
rect 1597 49 1601 53
rect 1580 38 1585 43
rect 1606 38 1611 43
rect 1584 28 1588 32
rect 1605 24 1609 28
rect 1597 12 1601 16
rect 1520 -3 1524 1
rect 1528 -12 1532 -8
rect 1596 -8 1600 -4
rect 1690 19 1694 23
rect 1663 13 1667 17
rect 1662 -7 1666 -3
rect 1705 -6 1709 -2
rect 1537 -44 1541 -40
rect 1596 -55 1600 -51
rect 1690 -18 1694 -14
rect 1727 -7 1731 -3
rect 1581 -68 1585 -64
rect 1605 -68 1609 -64
rect 1623 -86 1627 -82
rect 1596 -92 1600 -88
rect 1446 -116 1452 -110
rect 1447 -146 1453 -140
rect 1488 -147 1494 -141
rect 1401 -270 1405 -266
rect 1392 -290 1396 -286
rect 1322 -339 1326 -335
rect 1127 -355 1131 -351
rect 1067 -384 1071 -380
rect 1139 -385 1143 -381
rect 1082 -394 1086 -390
rect 1164 -385 1168 -381
rect 1186 -385 1190 -381
rect 1206 -377 1210 -373
rect 1216 -385 1220 -381
rect 1154 -395 1158 -391
rect 1240 -394 1244 -390
rect 1321 -370 1325 -366
rect 1273 -385 1277 -381
rect 1309 -382 1313 -378
rect 1272 -393 1276 -389
rect 1289 -390 1293 -386
rect 1299 -392 1303 -388
rect 1262 -400 1266 -396
rect 1348 -384 1352 -380
rect 1362 -391 1366 -387
rect 1331 -399 1335 -395
rect 1318 -409 1322 -405
rect 723 -432 728 -426
rect 407 -444 411 -440
rect 331 -480 336 -475
rect 379 -481 384 -476
rect 399 -492 403 -488
rect 509 -452 513 -447
rect 476 -464 480 -459
rect 472 -481 477 -476
rect 1009 -456 1013 -452
rect 565 -464 569 -460
rect 557 -481 562 -476
rect 323 -503 330 -496
rect 1369 -421 1373 -417
rect 1067 -431 1071 -427
rect 1105 -431 1109 -426
rect 1321 -428 1325 -424
rect 1158 -442 1162 -438
rect 1143 -452 1147 -448
rect 1244 -443 1248 -439
rect 1276 -444 1280 -440
rect 1168 -452 1172 -448
rect 1190 -452 1194 -448
rect 1220 -452 1224 -448
rect 1303 -445 1307 -441
rect 1277 -452 1281 -448
rect 1313 -455 1317 -451
rect 1210 -460 1214 -456
rect 1335 -438 1339 -434
rect 1366 -446 1370 -442
rect 1352 -453 1356 -449
rect 1322 -483 1326 -479
rect 1404 -360 1408 -356
rect 1404 -414 1408 -410
rect 1397 -445 1401 -441
rect 1546 -127 1550 -123
rect 1517 -236 1522 -230
rect 1467 -256 1471 -252
rect 1557 -134 1561 -130
rect 1690 -65 1694 -61
rect 1758 -61 1762 -57
rect 1766 -70 1770 -66
rect 1689 -85 1693 -81
rect 1689 -122 1693 -118
rect 1580 -144 1584 -140
rect 1606 -144 1610 -140
rect 1663 -130 1667 -126
rect 1739 -105 1745 -99
rect 1775 -106 1781 -100
rect 1691 -154 1695 -150
rect 1767 -153 1773 -147
rect 1623 -175 1627 -171
rect 1719 -177 1727 -169
rect 1598 -183 1602 -179
rect 1641 -186 1647 -180
rect 1666 -200 1672 -193
rect 1715 -203 1722 -195
rect 1765 -202 1771 -197
rect 1692 -222 1699 -216
rect 1642 -234 1647 -229
rect 1729 -231 1733 -227
rect 1758 -231 1762 -227
rect 1680 -246 1684 -242
rect 1557 -264 1561 -259
rect 1655 -254 1659 -250
rect 1727 -267 1734 -260
rect 1667 -285 1671 -281
rect 1698 -285 1702 -281
rect 1775 -277 1779 -273
rect 1737 -295 1741 -291
rect 1682 -337 1686 -333
rect 1655 -343 1659 -339
rect 1698 -364 1702 -360
rect 1682 -374 1686 -370
rect 1725 -338 1729 -334
rect 1718 -374 1722 -370
rect 1831 -310 1836 -304
rect 1452 -478 1460 -472
rect 1682 -421 1686 -417
rect 1734 -417 1738 -413
rect 1754 -417 1758 -413
rect 1681 -441 1685 -437
rect 1697 -452 1701 -448
rect 1721 -425 1725 -421
rect 1743 -425 1747 -421
rect 1681 -478 1685 -474
rect 1055 -494 1060 -489
rect 1655 -486 1659 -482
rect 1765 -443 1769 -439
rect 1740 -472 1744 -468
rect 1583 -505 1590 -498
rect 1607 -507 1612 -502
rect 1631 -507 1635 -502
rect 1306 -528 1313 -522
rect 1607 -528 1612 -522
rect 940 -540 949 -531
rect 1485 -541 1491 -534
rect 1013 -555 1020 -547
rect 1578 -558 1582 -554
rect 1355 -567 1360 -562
rect 1473 -566 1480 -558
rect 1683 -510 1687 -506
rect 1724 -501 1728 -497
rect 1653 -532 1658 -527
rect 1692 -532 1697 -527
rect 1654 -554 1659 -548
rect 1674 -555 1680 -550
rect 1693 -552 1697 -547
rect 1729 -558 1734 -553
rect 1640 -566 1645 -561
rect 1663 -576 1667 -572
rect 1755 -554 1759 -550
rect 1794 -568 1800 -562
rect 1806 -582 1813 -574
<< m3contact >>
rect 498 374 502 378
rect 517 353 521 357
rect 283 5 289 12
rect 1435 303 1440 308
rect 1515 280 1520 285
rect -12 -110 -8 -105
rect 525 -108 529 -104
rect 1300 38 1305 43
rect 1014 28 1019 33
rect 509 -132 513 -128
rect 528 -153 532 -149
rect 656 -189 660 -184
rect 687 -266 691 -262
rect 416 -373 421 -367
rect 952 -364 957 -360
rect 719 -404 724 -398
rect 687 -408 691 -404
rect 604 -430 609 -426
rect 909 -414 915 -408
rect 1301 -17 1305 -13
rect 1179 -26 1185 -19
rect 1501 -223 1507 -217
rect 1041 -336 1046 -332
rect 1501 -283 1506 -277
rect 626 -501 630 -497
rect 911 -538 916 -532
rect 1584 -545 1590 -539
rect 1602 -558 1606 -554
rect 1718 -557 1722 -553
rect 1823 -571 1830 -565
<< psubstratepcontact >>
rect 144 441 148 445
rect 231 441 235 445
rect 324 441 328 445
rect 536 443 540 447
rect 629 443 633 447
rect 716 443 720 447
rect 1571 439 1575 443
rect 1711 440 1715 444
rect 38 302 42 306
rect 116 302 120 306
rect 200 302 204 306
rect 270 302 274 306
rect 367 304 371 308
rect 445 304 449 308
rect 529 304 533 308
rect 1711 370 1715 374
rect 1571 361 1575 365
rect 599 304 603 308
rect 694 307 698 311
rect 772 307 776 311
rect 856 307 860 311
rect 1561 346 1565 350
rect 1721 329 1725 333
rect 1561 318 1565 322
rect 926 307 930 311
rect 131 292 135 296
rect 159 292 163 296
rect 460 294 464 298
rect 488 294 492 298
rect 787 297 791 301
rect 815 297 819 301
rect 1721 301 1725 305
rect 1711 286 1715 290
rect 1571 277 1575 281
rect 1378 242 1382 246
rect 1379 233 1383 237
rect 37 156 41 160
rect 115 156 119 160
rect 199 156 203 160
rect 269 156 273 160
rect 366 158 370 162
rect 444 158 448 162
rect 528 158 532 162
rect 1571 207 1575 211
rect 598 158 602 162
rect 693 161 697 165
rect 771 161 775 165
rect 855 161 859 165
rect 1711 208 1715 212
rect 925 161 929 165
rect 130 146 134 150
rect 158 146 162 150
rect 459 148 463 152
rect 487 148 491 152
rect 786 151 790 155
rect 814 151 818 155
rect 1378 102 1382 106
rect 1573 79 1577 83
rect 1713 80 1717 84
rect 331 8 335 12
rect 424 8 428 12
rect 511 8 515 12
rect 1713 10 1717 14
rect 1573 1 1577 5
rect 1563 -14 1567 -10
rect 1723 -31 1727 -27
rect 1563 -42 1567 -38
rect 155 -65 159 -61
rect 242 -65 246 -61
rect 335 -65 339 -61
rect 547 -63 551 -59
rect 640 -63 644 -59
rect 727 -63 731 -59
rect 1723 -59 1727 -55
rect 1713 -74 1717 -70
rect 1573 -83 1577 -79
rect 49 -204 53 -200
rect 127 -204 131 -200
rect 211 -204 215 -200
rect 281 -204 285 -200
rect 378 -202 382 -198
rect 456 -202 460 -198
rect 540 -202 544 -198
rect 1573 -153 1577 -149
rect 1713 -152 1717 -148
rect 610 -202 614 -198
rect 705 -199 709 -195
rect 783 -199 787 -195
rect 867 -199 871 -195
rect 937 -199 941 -195
rect 142 -214 146 -210
rect 170 -214 174 -210
rect 471 -212 475 -208
rect 499 -212 503 -208
rect 798 -209 802 -205
rect 826 -209 830 -205
rect 1410 -240 1414 -236
rect 48 -350 52 -346
rect 126 -350 130 -346
rect 210 -350 214 -346
rect 280 -350 284 -346
rect 377 -348 381 -344
rect 455 -348 459 -344
rect 539 -348 543 -344
rect 1705 -276 1709 -272
rect 609 -348 613 -344
rect 704 -345 708 -341
rect 782 -345 786 -341
rect 866 -345 870 -341
rect 936 -345 940 -341
rect 141 -360 145 -356
rect 169 -360 173 -356
rect 470 -358 474 -354
rect 498 -358 502 -354
rect 797 -355 801 -351
rect 825 -355 829 -351
rect 1705 -346 1709 -342
rect 1412 -393 1416 -389
rect 1715 -387 1719 -383
rect 1414 -419 1418 -415
rect 1715 -415 1719 -411
rect 1705 -430 1709 -426
rect 342 -498 346 -494
rect 435 -498 439 -494
rect 522 -498 526 -494
rect 1705 -508 1709 -504
<< nsubstratencontact >>
rect 1651 468 1655 472
rect 1651 454 1655 458
rect 1172 443 1176 447
rect 1226 443 1230 447
rect 1282 443 1286 447
rect 1336 443 1340 447
rect 1631 439 1635 443
rect 1651 440 1655 444
rect 1631 425 1635 429
rect 1631 411 1635 415
rect 1651 403 1655 407
rect 144 381 148 385
rect 231 381 235 385
rect 324 381 328 385
rect 536 383 540 387
rect 629 383 633 387
rect 716 383 720 387
rect 38 362 42 366
rect 52 362 56 366
rect 66 362 70 366
rect 149 362 153 366
rect 233 362 237 366
rect 270 362 274 366
rect 284 362 288 366
rect 298 362 302 366
rect 367 364 371 368
rect 381 364 385 368
rect 395 364 399 368
rect 478 364 482 368
rect 562 364 566 368
rect 599 364 603 368
rect 613 364 617 368
rect 627 364 631 368
rect 694 367 698 371
rect 708 367 712 371
rect 722 367 726 371
rect 805 367 809 371
rect 889 367 893 371
rect 926 367 930 371
rect 940 367 944 371
rect 954 367 958 371
rect 1176 316 1180 320
rect 1230 316 1234 320
rect 1286 316 1290 320
rect 1340 316 1344 320
rect 1501 318 1505 322
rect 1631 328 1635 332
rect 1651 319 1655 323
rect 1378 302 1382 306
rect 1172 298 1176 302
rect 1226 298 1230 302
rect 1282 298 1286 302
rect 1336 298 1340 302
rect 1781 329 1785 333
rect 159 232 163 236
rect 488 234 492 238
rect 815 237 819 241
rect 1631 244 1635 248
rect 37 216 41 220
rect 51 216 55 220
rect 65 216 69 220
rect 148 216 152 220
rect 232 216 236 220
rect 269 216 273 220
rect 283 216 287 220
rect 297 216 301 220
rect 366 218 370 222
rect 380 218 384 222
rect 394 218 398 222
rect 477 218 481 222
rect 561 218 565 222
rect 598 218 602 222
rect 612 218 616 222
rect 626 218 630 222
rect 693 221 697 225
rect 707 221 711 225
rect 721 221 725 225
rect 804 221 808 225
rect 888 221 892 225
rect 925 221 929 225
rect 939 221 943 225
rect 953 221 957 225
rect 1651 236 1655 240
rect 1651 222 1655 226
rect 1631 207 1635 211
rect 1651 208 1655 212
rect 1176 171 1180 175
rect 1230 171 1234 175
rect 1286 171 1290 175
rect 1340 171 1344 175
rect 1379 173 1383 177
rect 1631 193 1635 197
rect 1631 179 1635 183
rect 1378 162 1382 166
rect 1171 156 1175 160
rect 1225 156 1229 160
rect 1281 156 1285 160
rect 1335 156 1339 160
rect 1653 108 1657 112
rect 158 86 162 90
rect 487 88 491 92
rect 814 91 818 95
rect 1653 94 1657 98
rect 331 68 335 72
rect 424 68 428 72
rect 511 68 515 72
rect 1633 79 1637 83
rect 1653 80 1657 84
rect 1633 65 1637 69
rect 1633 51 1637 55
rect 1653 43 1657 47
rect 1175 29 1179 33
rect 1229 29 1233 33
rect 1285 29 1289 33
rect 1339 29 1343 33
rect 1503 -42 1507 -38
rect 1633 -32 1637 -28
rect 1653 -41 1657 -37
rect 1193 -68 1197 -64
rect 1247 -68 1251 -64
rect 1303 -68 1307 -64
rect 1357 -68 1361 -64
rect 1783 -31 1787 -27
rect 155 -125 159 -121
rect 242 -125 246 -121
rect 335 -125 339 -121
rect 547 -123 551 -119
rect 640 -123 644 -119
rect 727 -123 731 -119
rect 1633 -116 1637 -112
rect 1653 -124 1657 -120
rect 49 -144 53 -140
rect 63 -144 67 -140
rect 77 -144 81 -140
rect 160 -144 164 -140
rect 244 -144 248 -140
rect 281 -144 285 -140
rect 295 -144 299 -140
rect 309 -144 313 -140
rect 378 -142 382 -138
rect 392 -142 396 -138
rect 406 -142 410 -138
rect 489 -142 493 -138
rect 573 -142 577 -138
rect 610 -142 614 -138
rect 624 -142 628 -138
rect 638 -142 642 -138
rect 705 -139 709 -135
rect 719 -139 723 -135
rect 733 -139 737 -135
rect 816 -139 820 -135
rect 900 -139 904 -135
rect 937 -139 941 -135
rect 951 -139 955 -135
rect 965 -139 969 -135
rect 1653 -138 1657 -134
rect 1633 -153 1637 -149
rect 1653 -152 1657 -148
rect 1633 -167 1637 -163
rect 1633 -181 1637 -177
rect 1197 -195 1201 -191
rect 1251 -195 1255 -191
rect 1307 -195 1311 -191
rect 1361 -195 1365 -191
rect 1191 -213 1195 -209
rect 1245 -213 1249 -209
rect 1301 -213 1305 -209
rect 1355 -213 1359 -209
rect 170 -274 174 -270
rect 499 -272 503 -268
rect 826 -269 830 -265
rect 1645 -248 1649 -244
rect 1645 -262 1649 -258
rect 48 -290 52 -286
rect 62 -290 66 -286
rect 76 -290 80 -286
rect 159 -290 163 -286
rect 243 -290 247 -286
rect 280 -290 284 -286
rect 294 -290 298 -286
rect 308 -290 312 -286
rect 377 -288 381 -284
rect 391 -288 395 -284
rect 405 -288 409 -284
rect 488 -288 492 -284
rect 572 -288 576 -284
rect 609 -288 613 -284
rect 623 -288 627 -284
rect 637 -288 641 -284
rect 704 -285 708 -281
rect 718 -285 722 -281
rect 732 -285 736 -281
rect 815 -285 819 -281
rect 899 -285 903 -281
rect 936 -285 940 -281
rect 950 -285 954 -281
rect 964 -285 968 -281
rect 1410 -300 1414 -296
rect 1645 -276 1649 -272
rect 1645 -313 1649 -309
rect 1412 -333 1416 -329
rect 1195 -340 1199 -336
rect 1249 -340 1253 -336
rect 1305 -340 1309 -336
rect 1359 -340 1363 -336
rect 1192 -355 1196 -351
rect 1246 -355 1250 -351
rect 1302 -355 1306 -351
rect 1356 -355 1360 -351
rect 1645 -397 1649 -393
rect 169 -420 173 -416
rect 498 -418 502 -414
rect 825 -415 829 -411
rect 342 -438 346 -434
rect 435 -438 439 -434
rect 522 -438 526 -434
rect 1775 -387 1779 -383
rect 1196 -482 1200 -478
rect 1250 -482 1254 -478
rect 1306 -482 1310 -478
rect 1360 -482 1364 -478
rect 1414 -479 1418 -475
rect 1645 -480 1649 -476
rect 1645 -494 1649 -490
rect 1645 -508 1649 -504
<< psubstratepdiff >>
rect 535 447 541 448
rect 143 445 149 446
rect 143 441 144 445
rect 148 441 149 445
rect 143 440 149 441
rect 230 445 236 446
rect 230 441 231 445
rect 235 441 236 445
rect 230 440 236 441
rect 323 445 329 446
rect 323 441 324 445
rect 328 441 329 445
rect 535 443 536 447
rect 540 443 541 447
rect 535 442 541 443
rect 628 447 634 448
rect 628 443 629 447
rect 633 443 634 447
rect 323 440 329 441
rect 628 442 634 443
rect 715 447 721 448
rect 715 443 716 447
rect 720 443 721 447
rect 715 442 721 443
rect 1570 443 1576 444
rect 1570 439 1571 443
rect 1575 439 1576 443
rect 1570 438 1576 439
rect 1710 444 1716 445
rect 1710 440 1711 444
rect 1715 440 1716 444
rect 1710 439 1716 440
rect 37 306 43 307
rect 37 302 38 306
rect 42 302 43 306
rect 37 301 43 302
rect 115 306 121 307
rect 115 302 116 306
rect 120 302 121 306
rect 115 301 121 302
rect 199 306 205 307
rect 199 302 200 306
rect 204 302 205 306
rect 199 301 205 302
rect 366 308 372 309
rect 269 306 275 307
rect 269 302 270 306
rect 274 302 275 306
rect 269 301 275 302
rect 366 304 367 308
rect 371 304 372 308
rect 366 303 372 304
rect 444 308 450 309
rect 444 304 445 308
rect 449 304 450 308
rect 444 303 450 304
rect 528 308 534 309
rect 528 304 529 308
rect 533 304 534 308
rect 528 303 534 304
rect 1710 374 1716 375
rect 1710 370 1711 374
rect 1715 370 1716 374
rect 1710 369 1716 370
rect 1570 365 1576 366
rect 1570 361 1571 365
rect 1575 361 1576 365
rect 1570 360 1576 361
rect 693 311 699 312
rect 598 308 604 309
rect 598 304 599 308
rect 603 304 604 308
rect 598 303 604 304
rect 693 307 694 311
rect 698 307 699 311
rect 693 306 699 307
rect 771 311 777 312
rect 771 307 772 311
rect 776 307 777 311
rect 771 306 777 307
rect 855 311 861 312
rect 855 307 856 311
rect 860 307 861 311
rect 855 306 861 307
rect 1560 350 1566 351
rect 1560 346 1561 350
rect 1565 346 1566 350
rect 1560 322 1566 346
rect 1720 333 1726 334
rect 1720 329 1721 333
rect 1725 329 1726 333
rect 1560 318 1561 322
rect 1565 318 1566 322
rect 1560 317 1566 318
rect 925 311 931 312
rect 925 307 926 311
rect 930 307 931 311
rect 925 306 931 307
rect 786 301 820 302
rect 459 298 493 299
rect 130 296 164 297
rect 130 292 131 296
rect 135 292 159 296
rect 163 292 164 296
rect 459 294 460 298
rect 464 294 488 298
rect 492 294 493 298
rect 786 297 787 301
rect 791 297 815 301
rect 819 297 820 301
rect 786 296 820 297
rect 459 293 493 294
rect 130 291 164 292
rect 1720 305 1726 329
rect 1720 301 1721 305
rect 1725 301 1726 305
rect 1720 300 1726 301
rect 1710 290 1716 291
rect 1710 286 1711 290
rect 1715 286 1716 290
rect 1710 285 1716 286
rect 1570 281 1576 282
rect 1570 277 1571 281
rect 1575 277 1576 281
rect 1570 276 1576 277
rect 1377 246 1383 247
rect 1377 242 1378 246
rect 1382 242 1383 246
rect 1377 241 1383 242
rect 1378 237 1384 238
rect 1378 233 1379 237
rect 1383 233 1384 237
rect 1378 232 1384 233
rect 36 160 42 161
rect 36 156 37 160
rect 41 156 42 160
rect 36 155 42 156
rect 114 160 120 161
rect 114 156 115 160
rect 119 156 120 160
rect 114 155 120 156
rect 198 160 204 161
rect 198 156 199 160
rect 203 156 204 160
rect 198 155 204 156
rect 365 162 371 163
rect 268 160 274 161
rect 268 156 269 160
rect 273 156 274 160
rect 268 155 274 156
rect 365 158 366 162
rect 370 158 371 162
rect 365 157 371 158
rect 443 162 449 163
rect 443 158 444 162
rect 448 158 449 162
rect 443 157 449 158
rect 527 162 533 163
rect 527 158 528 162
rect 532 158 533 162
rect 527 157 533 158
rect 1570 211 1576 212
rect 1570 207 1571 211
rect 1575 207 1576 211
rect 1570 206 1576 207
rect 692 165 698 166
rect 597 162 603 163
rect 597 158 598 162
rect 602 158 603 162
rect 597 157 603 158
rect 692 161 693 165
rect 697 161 698 165
rect 692 160 698 161
rect 770 165 776 166
rect 770 161 771 165
rect 775 161 776 165
rect 770 160 776 161
rect 854 165 860 166
rect 854 161 855 165
rect 859 161 860 165
rect 854 160 860 161
rect 1710 212 1716 213
rect 1710 208 1711 212
rect 1715 208 1716 212
rect 1710 207 1716 208
rect 924 165 930 166
rect 924 161 925 165
rect 929 161 930 165
rect 924 160 930 161
rect 785 155 819 156
rect 458 152 492 153
rect 129 150 163 151
rect 129 146 130 150
rect 134 146 158 150
rect 162 146 163 150
rect 458 148 459 152
rect 463 148 487 152
rect 491 148 492 152
rect 785 151 786 155
rect 790 151 814 155
rect 818 151 819 155
rect 785 150 819 151
rect 458 147 492 148
rect 129 145 163 146
rect 1377 106 1383 107
rect 1377 102 1378 106
rect 1382 102 1383 106
rect 1377 101 1383 102
rect 1572 83 1578 84
rect 1572 79 1573 83
rect 1577 79 1578 83
rect 1572 78 1578 79
rect 1712 84 1718 85
rect 1712 80 1713 84
rect 1717 80 1718 84
rect 1712 79 1718 80
rect 330 12 336 13
rect 330 8 331 12
rect 335 8 336 12
rect 330 7 336 8
rect 423 12 429 13
rect 423 8 424 12
rect 428 8 429 12
rect 423 7 429 8
rect 510 12 516 13
rect 510 8 511 12
rect 515 8 516 12
rect 510 7 516 8
rect 1712 14 1718 15
rect 1712 10 1713 14
rect 1717 10 1718 14
rect 1712 9 1718 10
rect 1572 5 1578 6
rect 1572 1 1573 5
rect 1577 1 1578 5
rect 1572 0 1578 1
rect 1562 -10 1568 -9
rect 1562 -14 1563 -10
rect 1567 -14 1568 -10
rect 1562 -38 1568 -14
rect 1722 -27 1728 -26
rect 1722 -31 1723 -27
rect 1727 -31 1728 -27
rect 1562 -42 1563 -38
rect 1567 -42 1568 -38
rect 1562 -43 1568 -42
rect 546 -59 552 -58
rect 154 -61 160 -60
rect 154 -65 155 -61
rect 159 -65 160 -61
rect 154 -66 160 -65
rect 241 -61 247 -60
rect 241 -65 242 -61
rect 246 -65 247 -61
rect 241 -66 247 -65
rect 334 -61 340 -60
rect 334 -65 335 -61
rect 339 -65 340 -61
rect 546 -63 547 -59
rect 551 -63 552 -59
rect 546 -64 552 -63
rect 639 -59 645 -58
rect 639 -63 640 -59
rect 644 -63 645 -59
rect 334 -66 340 -65
rect 639 -64 645 -63
rect 726 -59 732 -58
rect 726 -63 727 -59
rect 731 -63 732 -59
rect 726 -64 732 -63
rect 1722 -55 1728 -31
rect 1722 -59 1723 -55
rect 1727 -59 1728 -55
rect 1722 -60 1728 -59
rect 1712 -70 1718 -69
rect 1712 -74 1713 -70
rect 1717 -74 1718 -70
rect 1712 -75 1718 -74
rect 1572 -79 1578 -78
rect 1572 -83 1573 -79
rect 1577 -83 1578 -79
rect 1572 -84 1578 -83
rect 48 -200 54 -199
rect 48 -204 49 -200
rect 53 -204 54 -200
rect 48 -205 54 -204
rect 126 -200 132 -199
rect 126 -204 127 -200
rect 131 -204 132 -200
rect 126 -205 132 -204
rect 210 -200 216 -199
rect 210 -204 211 -200
rect 215 -204 216 -200
rect 210 -205 216 -204
rect 377 -198 383 -197
rect 280 -200 286 -199
rect 280 -204 281 -200
rect 285 -204 286 -200
rect 280 -205 286 -204
rect 377 -202 378 -198
rect 382 -202 383 -198
rect 377 -203 383 -202
rect 455 -198 461 -197
rect 455 -202 456 -198
rect 460 -202 461 -198
rect 455 -203 461 -202
rect 539 -198 545 -197
rect 539 -202 540 -198
rect 544 -202 545 -198
rect 539 -203 545 -202
rect 1572 -149 1578 -148
rect 1572 -153 1573 -149
rect 1577 -153 1578 -149
rect 1572 -154 1578 -153
rect 1712 -148 1718 -147
rect 1712 -152 1713 -148
rect 1717 -152 1718 -148
rect 1712 -153 1718 -152
rect 704 -195 710 -194
rect 609 -198 615 -197
rect 609 -202 610 -198
rect 614 -202 615 -198
rect 609 -203 615 -202
rect 704 -199 705 -195
rect 709 -199 710 -195
rect 704 -200 710 -199
rect 782 -195 788 -194
rect 782 -199 783 -195
rect 787 -199 788 -195
rect 782 -200 788 -199
rect 866 -195 872 -194
rect 866 -199 867 -195
rect 871 -199 872 -195
rect 866 -200 872 -199
rect 936 -195 942 -194
rect 936 -199 937 -195
rect 941 -199 942 -195
rect 936 -200 942 -199
rect 797 -205 831 -204
rect 470 -208 504 -207
rect 141 -210 175 -209
rect 141 -214 142 -210
rect 146 -214 170 -210
rect 174 -214 175 -210
rect 470 -212 471 -208
rect 475 -212 499 -208
rect 503 -212 504 -208
rect 797 -209 798 -205
rect 802 -209 826 -205
rect 830 -209 831 -205
rect 797 -210 831 -209
rect 470 -213 504 -212
rect 141 -215 175 -214
rect 1409 -236 1415 -235
rect 1409 -240 1410 -236
rect 1414 -240 1415 -236
rect 1409 -241 1415 -240
rect 47 -346 53 -345
rect 47 -350 48 -346
rect 52 -350 53 -346
rect 47 -351 53 -350
rect 125 -346 131 -345
rect 125 -350 126 -346
rect 130 -350 131 -346
rect 125 -351 131 -350
rect 209 -346 215 -345
rect 209 -350 210 -346
rect 214 -350 215 -346
rect 209 -351 215 -350
rect 376 -344 382 -343
rect 279 -346 285 -345
rect 279 -350 280 -346
rect 284 -350 285 -346
rect 279 -351 285 -350
rect 376 -348 377 -344
rect 381 -348 382 -344
rect 376 -349 382 -348
rect 454 -344 460 -343
rect 454 -348 455 -344
rect 459 -348 460 -344
rect 454 -349 460 -348
rect 538 -344 544 -343
rect 538 -348 539 -344
rect 543 -348 544 -344
rect 538 -349 544 -348
rect 1704 -272 1710 -271
rect 1704 -276 1705 -272
rect 1709 -276 1710 -272
rect 1704 -277 1710 -276
rect 703 -341 709 -340
rect 608 -344 614 -343
rect 608 -348 609 -344
rect 613 -348 614 -344
rect 608 -349 614 -348
rect 703 -345 704 -341
rect 708 -345 709 -341
rect 703 -346 709 -345
rect 781 -341 787 -340
rect 781 -345 782 -341
rect 786 -345 787 -341
rect 781 -346 787 -345
rect 865 -341 871 -340
rect 865 -345 866 -341
rect 870 -345 871 -341
rect 865 -346 871 -345
rect 935 -341 941 -340
rect 935 -345 936 -341
rect 940 -345 941 -341
rect 935 -346 941 -345
rect 796 -351 830 -350
rect 469 -354 503 -353
rect 140 -356 174 -355
rect 140 -360 141 -356
rect 145 -360 169 -356
rect 173 -360 174 -356
rect 469 -358 470 -354
rect 474 -358 498 -354
rect 502 -358 503 -354
rect 796 -355 797 -351
rect 801 -355 825 -351
rect 829 -355 830 -351
rect 796 -356 830 -355
rect 469 -359 503 -358
rect 140 -361 174 -360
rect 1704 -342 1710 -341
rect 1704 -346 1705 -342
rect 1709 -346 1710 -342
rect 1704 -347 1710 -346
rect 1411 -389 1417 -388
rect 1411 -393 1412 -389
rect 1416 -393 1417 -389
rect 1714 -383 1720 -382
rect 1714 -387 1715 -383
rect 1719 -387 1720 -383
rect 1411 -394 1417 -393
rect 1413 -415 1419 -414
rect 1413 -419 1414 -415
rect 1418 -419 1419 -415
rect 1413 -420 1419 -419
rect 1714 -411 1720 -387
rect 1714 -415 1715 -411
rect 1719 -415 1720 -411
rect 1714 -416 1720 -415
rect 1704 -426 1710 -425
rect 1704 -430 1705 -426
rect 1709 -430 1710 -426
rect 1704 -431 1710 -430
rect 341 -494 347 -493
rect 341 -498 342 -494
rect 346 -498 347 -494
rect 341 -499 347 -498
rect 434 -494 440 -493
rect 434 -498 435 -494
rect 439 -498 440 -494
rect 434 -499 440 -498
rect 521 -494 527 -493
rect 521 -498 522 -494
rect 526 -498 527 -494
rect 521 -499 527 -498
rect 1704 -504 1710 -503
rect 1704 -508 1705 -504
rect 1709 -508 1710 -504
rect 1704 -509 1710 -508
<< nsubstratendiff >>
rect 1650 472 1656 473
rect 1650 468 1651 472
rect 1655 468 1656 472
rect 1650 458 1656 468
rect 1650 454 1651 458
rect 1655 454 1656 458
rect 1650 444 1656 454
rect 1630 443 1636 444
rect 1630 439 1631 443
rect 1635 439 1636 443
rect 1650 440 1651 444
rect 1655 440 1656 444
rect 1650 439 1656 440
rect 1630 429 1636 439
rect 143 385 149 386
rect 230 385 236 386
rect 535 387 541 388
rect 1630 425 1631 429
rect 1635 425 1636 429
rect 628 387 634 388
rect 715 387 721 388
rect 1630 415 1636 425
rect 1630 411 1631 415
rect 1635 411 1636 415
rect 1630 410 1636 411
rect 1650 407 1656 408
rect 1650 403 1651 407
rect 1655 403 1656 407
rect 1650 402 1656 403
rect 323 385 329 386
rect 143 381 144 385
rect 148 381 149 385
rect 143 380 149 381
rect 230 381 231 385
rect 235 381 236 385
rect 230 380 236 381
rect 323 381 324 385
rect 328 381 329 385
rect 535 383 536 387
rect 540 383 541 387
rect 535 382 541 383
rect 628 383 629 387
rect 633 383 634 387
rect 628 382 634 383
rect 715 383 716 387
rect 720 383 721 387
rect 715 382 721 383
rect 323 380 329 381
rect 366 368 400 369
rect 37 366 71 367
rect 37 362 38 366
rect 42 362 52 366
rect 56 362 66 366
rect 70 362 71 366
rect 148 366 154 367
rect 37 361 71 362
rect 148 362 149 366
rect 153 362 154 366
rect 232 366 238 367
rect 148 361 154 362
rect 232 362 233 366
rect 237 362 238 366
rect 269 366 303 367
rect 232 361 238 362
rect 269 362 270 366
rect 274 362 284 366
rect 288 362 298 366
rect 302 362 303 366
rect 366 364 367 368
rect 371 364 381 368
rect 385 364 395 368
rect 399 364 400 368
rect 477 368 483 369
rect 366 363 400 364
rect 269 361 303 362
rect 477 364 478 368
rect 482 364 483 368
rect 561 368 567 369
rect 477 363 483 364
rect 561 364 562 368
rect 566 364 567 368
rect 598 368 632 369
rect 561 363 567 364
rect 598 364 599 368
rect 603 364 613 368
rect 617 364 627 368
rect 631 364 632 368
rect 693 367 694 371
rect 698 367 708 371
rect 712 367 722 371
rect 726 367 727 371
rect 804 371 810 372
rect 693 366 727 367
rect 598 363 632 364
rect 804 367 805 371
rect 809 367 810 371
rect 888 371 894 372
rect 804 366 810 367
rect 888 367 889 371
rect 893 367 894 371
rect 925 371 959 372
rect 888 366 894 367
rect 925 367 926 371
rect 930 367 940 371
rect 944 367 954 371
rect 958 367 959 371
rect 925 366 959 367
rect 1500 322 1506 323
rect 1500 318 1501 322
rect 1505 318 1506 322
rect 1500 317 1506 318
rect 1630 332 1636 333
rect 1630 328 1631 332
rect 1635 328 1636 332
rect 1630 327 1636 328
rect 1650 323 1656 324
rect 1650 319 1651 323
rect 1655 319 1656 323
rect 1650 318 1656 319
rect 1377 306 1383 307
rect 1377 302 1378 306
rect 1382 302 1383 306
rect 1377 301 1383 302
rect 1780 333 1786 334
rect 1780 329 1781 333
rect 1785 329 1786 333
rect 1780 328 1786 329
rect 158 236 164 237
rect 814 241 820 242
rect 487 238 493 239
rect 158 232 159 236
rect 163 232 164 236
rect 487 234 488 238
rect 492 234 493 238
rect 814 237 815 241
rect 819 237 820 241
rect 1630 248 1636 249
rect 1630 244 1631 248
rect 1635 244 1636 248
rect 1630 243 1636 244
rect 1650 240 1656 241
rect 814 236 820 237
rect 487 233 493 234
rect 158 231 164 232
rect 692 225 726 226
rect 365 222 399 223
rect 36 220 70 221
rect 36 216 37 220
rect 41 216 51 220
rect 55 216 65 220
rect 69 216 70 220
rect 147 220 153 221
rect 36 215 70 216
rect 147 216 148 220
rect 152 216 153 220
rect 231 220 237 221
rect 147 215 153 216
rect 231 216 232 220
rect 236 216 237 220
rect 268 220 302 221
rect 231 215 237 216
rect 268 216 269 220
rect 273 216 283 220
rect 287 216 297 220
rect 301 216 302 220
rect 365 218 366 222
rect 370 218 380 222
rect 384 218 394 222
rect 398 218 399 222
rect 476 222 482 223
rect 365 217 399 218
rect 268 215 302 216
rect 476 218 477 222
rect 481 218 482 222
rect 560 222 566 223
rect 476 217 482 218
rect 560 218 561 222
rect 565 218 566 222
rect 597 222 631 223
rect 560 217 566 218
rect 597 218 598 222
rect 602 218 612 222
rect 616 218 626 222
rect 630 218 631 222
rect 692 221 693 225
rect 697 221 707 225
rect 711 221 721 225
rect 725 221 726 225
rect 803 225 809 226
rect 692 220 726 221
rect 597 217 631 218
rect 803 221 804 225
rect 808 221 809 225
rect 887 225 893 226
rect 803 220 809 221
rect 887 221 888 225
rect 892 221 893 225
rect 924 225 958 226
rect 887 220 893 221
rect 924 221 925 225
rect 929 221 939 225
rect 943 221 953 225
rect 957 221 958 225
rect 924 220 958 221
rect 1650 236 1651 240
rect 1655 236 1656 240
rect 1650 226 1656 236
rect 1650 222 1651 226
rect 1655 222 1656 226
rect 1650 212 1656 222
rect 1630 211 1636 212
rect 1630 207 1631 211
rect 1635 207 1636 211
rect 1650 208 1651 212
rect 1655 208 1656 212
rect 1650 207 1656 208
rect 1378 177 1384 178
rect 1378 173 1379 177
rect 1383 173 1384 177
rect 1378 172 1384 173
rect 1630 197 1636 207
rect 1630 193 1631 197
rect 1635 193 1636 197
rect 1630 183 1636 193
rect 1630 179 1631 183
rect 1635 179 1636 183
rect 1630 178 1636 179
rect 1377 166 1383 167
rect 1377 162 1378 166
rect 1382 162 1383 166
rect 1377 161 1383 162
rect 157 90 163 91
rect 1652 112 1658 113
rect 1652 108 1653 112
rect 1657 108 1658 112
rect 1652 98 1658 108
rect 813 95 819 96
rect 486 92 492 93
rect 157 86 158 90
rect 162 86 163 90
rect 486 88 487 92
rect 491 88 492 92
rect 813 91 814 95
rect 818 91 819 95
rect 813 90 819 91
rect 1652 94 1653 98
rect 1657 94 1658 98
rect 486 87 492 88
rect 157 85 163 86
rect 330 72 336 73
rect 330 68 331 72
rect 335 68 336 72
rect 423 72 429 73
rect 423 68 424 72
rect 428 68 429 72
rect 510 72 516 73
rect 510 68 511 72
rect 515 68 516 72
rect 330 67 336 68
rect 423 67 429 68
rect 510 67 516 68
rect 1652 84 1658 94
rect 1632 83 1638 84
rect 1632 79 1633 83
rect 1637 79 1638 83
rect 1652 80 1653 84
rect 1657 80 1658 84
rect 1652 79 1658 80
rect 1632 69 1638 79
rect 1632 65 1633 69
rect 1637 65 1638 69
rect 1632 55 1638 65
rect 1632 51 1633 55
rect 1637 51 1638 55
rect 1632 50 1638 51
rect 1652 47 1658 48
rect 1652 43 1653 47
rect 1657 43 1658 47
rect 1652 42 1658 43
rect 1502 -38 1508 -37
rect 1502 -42 1503 -38
rect 1507 -42 1508 -38
rect 1502 -43 1508 -42
rect 1632 -28 1638 -27
rect 1632 -32 1633 -28
rect 1637 -32 1638 -28
rect 1632 -33 1638 -32
rect 1652 -37 1658 -36
rect 1652 -41 1653 -37
rect 1657 -41 1658 -37
rect 1652 -42 1658 -41
rect 1782 -27 1788 -26
rect 1782 -31 1783 -27
rect 1787 -31 1788 -27
rect 1782 -32 1788 -31
rect 154 -121 160 -120
rect 241 -121 247 -120
rect 546 -119 552 -118
rect 639 -119 645 -118
rect 726 -119 732 -118
rect 334 -121 340 -120
rect 154 -125 155 -121
rect 159 -125 160 -121
rect 154 -126 160 -125
rect 241 -125 242 -121
rect 246 -125 247 -121
rect 241 -126 247 -125
rect 334 -125 335 -121
rect 339 -125 340 -121
rect 546 -123 547 -119
rect 551 -123 552 -119
rect 546 -124 552 -123
rect 639 -123 640 -119
rect 644 -123 645 -119
rect 639 -124 645 -123
rect 726 -123 727 -119
rect 731 -123 732 -119
rect 1632 -112 1638 -111
rect 1632 -116 1633 -112
rect 1637 -116 1638 -112
rect 1632 -117 1638 -116
rect 1652 -120 1658 -119
rect 726 -124 732 -123
rect 334 -126 340 -125
rect 1652 -124 1653 -120
rect 1657 -124 1658 -120
rect 377 -138 411 -137
rect 48 -140 82 -139
rect 48 -144 49 -140
rect 53 -144 63 -140
rect 67 -144 77 -140
rect 81 -144 82 -140
rect 159 -140 165 -139
rect 48 -145 82 -144
rect 159 -144 160 -140
rect 164 -144 165 -140
rect 243 -140 249 -139
rect 159 -145 165 -144
rect 243 -144 244 -140
rect 248 -144 249 -140
rect 280 -140 314 -139
rect 243 -145 249 -144
rect 280 -144 281 -140
rect 285 -144 295 -140
rect 299 -144 309 -140
rect 313 -144 314 -140
rect 377 -142 378 -138
rect 382 -142 392 -138
rect 396 -142 406 -138
rect 410 -142 411 -138
rect 488 -138 494 -137
rect 377 -143 411 -142
rect 280 -145 314 -144
rect 488 -142 489 -138
rect 493 -142 494 -138
rect 572 -138 578 -137
rect 488 -143 494 -142
rect 572 -142 573 -138
rect 577 -142 578 -138
rect 609 -138 643 -137
rect 572 -143 578 -142
rect 609 -142 610 -138
rect 614 -142 624 -138
rect 628 -142 638 -138
rect 642 -142 643 -138
rect 704 -139 705 -135
rect 709 -139 719 -135
rect 723 -139 733 -135
rect 737 -139 738 -135
rect 815 -135 821 -134
rect 704 -140 738 -139
rect 609 -143 643 -142
rect 815 -139 816 -135
rect 820 -139 821 -135
rect 899 -135 905 -134
rect 815 -140 821 -139
rect 899 -139 900 -135
rect 904 -139 905 -135
rect 936 -135 970 -134
rect 899 -140 905 -139
rect 936 -139 937 -135
rect 941 -139 951 -135
rect 955 -139 965 -135
rect 969 -139 970 -135
rect 1652 -134 1658 -124
rect 1652 -138 1653 -134
rect 1657 -138 1658 -134
rect 936 -140 970 -139
rect 1652 -148 1658 -138
rect 1632 -149 1638 -148
rect 1632 -153 1633 -149
rect 1637 -153 1638 -149
rect 1652 -152 1653 -148
rect 1657 -152 1658 -148
rect 1652 -153 1658 -152
rect 1632 -163 1638 -153
rect 1632 -167 1633 -163
rect 1637 -167 1638 -163
rect 1632 -177 1638 -167
rect 1632 -181 1633 -177
rect 1637 -181 1638 -177
rect 1632 -182 1638 -181
rect 169 -270 175 -269
rect 825 -265 831 -264
rect 498 -268 504 -267
rect 169 -274 170 -270
rect 174 -274 175 -270
rect 498 -272 499 -268
rect 503 -272 504 -268
rect 825 -269 826 -265
rect 830 -269 831 -265
rect 1644 -244 1650 -243
rect 1644 -248 1645 -244
rect 1649 -248 1650 -244
rect 1644 -258 1650 -248
rect 825 -270 831 -269
rect 1644 -262 1645 -258
rect 1649 -262 1650 -258
rect 498 -273 504 -272
rect 169 -275 175 -274
rect 703 -281 737 -280
rect 376 -284 410 -283
rect 47 -286 81 -285
rect 47 -290 48 -286
rect 52 -290 62 -286
rect 66 -290 76 -286
rect 80 -290 81 -286
rect 158 -286 164 -285
rect 47 -291 81 -290
rect 158 -290 159 -286
rect 163 -290 164 -286
rect 242 -286 248 -285
rect 158 -291 164 -290
rect 242 -290 243 -286
rect 247 -290 248 -286
rect 279 -286 313 -285
rect 242 -291 248 -290
rect 279 -290 280 -286
rect 284 -290 294 -286
rect 298 -290 308 -286
rect 312 -290 313 -286
rect 376 -288 377 -284
rect 381 -288 391 -284
rect 395 -288 405 -284
rect 409 -288 410 -284
rect 487 -284 493 -283
rect 376 -289 410 -288
rect 279 -291 313 -290
rect 487 -288 488 -284
rect 492 -288 493 -284
rect 571 -284 577 -283
rect 487 -289 493 -288
rect 571 -288 572 -284
rect 576 -288 577 -284
rect 608 -284 642 -283
rect 571 -289 577 -288
rect 608 -288 609 -284
rect 613 -288 623 -284
rect 627 -288 637 -284
rect 641 -288 642 -284
rect 703 -285 704 -281
rect 708 -285 718 -281
rect 722 -285 732 -281
rect 736 -285 737 -281
rect 814 -281 820 -280
rect 703 -286 737 -285
rect 608 -289 642 -288
rect 814 -285 815 -281
rect 819 -285 820 -281
rect 898 -281 904 -280
rect 814 -286 820 -285
rect 898 -285 899 -281
rect 903 -285 904 -281
rect 935 -281 969 -280
rect 898 -286 904 -285
rect 935 -285 936 -281
rect 940 -285 950 -281
rect 954 -285 964 -281
rect 968 -285 969 -281
rect 935 -286 969 -285
rect 1409 -296 1415 -295
rect 1409 -300 1410 -296
rect 1414 -300 1415 -296
rect 1409 -301 1415 -300
rect 1644 -272 1650 -262
rect 1644 -276 1645 -272
rect 1649 -276 1650 -272
rect 1644 -277 1650 -276
rect 1644 -309 1650 -308
rect 1644 -313 1645 -309
rect 1649 -313 1650 -309
rect 1644 -314 1650 -313
rect 1411 -329 1417 -328
rect 1411 -333 1412 -329
rect 1416 -333 1417 -329
rect 1411 -334 1417 -333
rect 168 -416 174 -415
rect 1644 -393 1650 -392
rect 1644 -397 1645 -393
rect 1649 -397 1650 -393
rect 1644 -398 1650 -397
rect 824 -411 830 -410
rect 497 -414 503 -413
rect 168 -420 169 -416
rect 173 -420 174 -416
rect 497 -418 498 -414
rect 502 -418 503 -414
rect 824 -415 825 -411
rect 829 -415 830 -411
rect 824 -416 830 -415
rect 497 -419 503 -418
rect 168 -421 174 -420
rect 341 -434 347 -433
rect 341 -438 342 -434
rect 346 -438 347 -434
rect 434 -434 440 -433
rect 434 -438 435 -434
rect 439 -438 440 -434
rect 521 -434 527 -433
rect 521 -438 522 -434
rect 526 -438 527 -434
rect 341 -439 347 -438
rect 434 -439 440 -438
rect 521 -439 527 -438
rect 1774 -383 1780 -382
rect 1774 -387 1775 -383
rect 1779 -387 1780 -383
rect 1774 -388 1780 -387
rect 1413 -475 1419 -474
rect 1413 -479 1414 -475
rect 1418 -479 1419 -475
rect 1413 -480 1419 -479
rect 1644 -476 1650 -475
rect 1644 -480 1645 -476
rect 1649 -480 1650 -476
rect 1644 -490 1650 -480
rect 1644 -494 1645 -490
rect 1649 -494 1650 -490
rect 1644 -504 1650 -494
rect 1644 -508 1645 -504
rect 1649 -508 1650 -504
rect 1644 -509 1650 -508
<< pad >>
rect 171 375 175 379
rect 182 -131 186 -127
<< labels >>
rlabel metal1 802 91 802 91 2 vdd
rlabel m2contact 112 425 112 425 1 q0_M1
rlabel metal1 148 417 148 417 1 q0b2_M1
rlabel metal1 320 424 320 424 1 q0b0_n_M1
rlabel metal1 440 430 440 430 1 b2_M1
rlabel metal1 441 409 441 409 1 b1_M1
rlabel metal1 441 390 441 390 1 b0_M1
rlabel metal1 535 428 535 428 1 q1b0_M1
rlabel metal1 637 435 637 435 1 q1b1_M1
rlabel metal1 637 413 637 413 1 q1b1_n_M1
rlabel metal1 715 424 715 424 1 q1b2_M1
rlabel metal1 724 424 724 424 1 q1b2_n_M1
rlabel m2contact 751 427 751 427 1 q1_M1
rlabel metal1 940 335 940 335 1 zc1_n_3_M1
rlabel metal1 926 335 926 335 1 c1_3_M1
rlabel metal1 912 339 912 339 1 s_fa3_M1
rlabel metal1 889 357 889 357 1 cn_3_M1
rlabel metal1 828 339 828 339 1 so_3_M1
rlabel metal1 816 360 816 360 1 bn3_M1
rlabel ptransistor 812 344 812 344 1 an3_M1
rlabel metal1 715 339 715 339 1 co_n3_M1
rlabel metal1 702 319 702 319 1 co_3_M1
rlabel metal1 599 332 599 332 1 c1_2_M1
rlabel metal1 613 332 613 332 1 zc1_2_n_M1
rlabel ntransistor 578 319 578 319 1 son_2_M1
rlabel pdcontact 575 349 575 349 1 s_fa2_M1
rlabel metal1 563 332 563 332 1 cn2_M1
rlabel metal1 501 336 501 336 1 so_2_M1
rlabel polycontact 491 332 491 332 1 an_2_M1
rlabel polycontact 485 333 485 333 1 bn_2_M1
rlabel metal1 388 335 388 335 1 co_n2_M1
rlabel metal1 375 316 375 316 1 co_2_M1
rlabel metal1 284 330 284 330 1 zc1_n1_M1
rlabel metal1 270 330 270 330 1 c1_1_M1
rlabel ntransistor 249 317 249 317 1 a1_n_M1
rlabel ntransistor 165 318 165 318 1 an_1_M1
rlabel metal1 172 334 172 334 1 so_1_M1
rlabel metal1 59 334 59 334 1 co_n1_M1
rlabel metal1 46 314 46 314 1 co_1_M1
rlabel metal1 155 262 155 262 1 c_fa1_n_M1
rlabel metal1 163 262 163 262 1 c_fa1_M1
rlabel metal1 484 266 484 266 1 c_fa_n_M1
rlabel metal1 492 270 492 270 1 c_fa2_M1
rlabel metal1 811 269 811 269 1 c_fa3_n_M1
rlabel metal1 819 273 819 273 1 c_fa3_M1
rlabel metal1 939 189 939 189 1 zc1_6_n_M1
rlabel metal1 925 189 925 189 1 c1_6_M1
rlabel ntransistor 904 176 904 176 1 s_fa_6_n_M1
rlabel metal1 887 210 887 210 1 cn_6_M1
rlabel metal1 827 193 827 193 1 so_6_M1
rlabel ptransistor 811 198 811 198 1 an_6_M1
rlabel metal1 772 187 772 187 1 bn_6_M1
rlabel metal1 714 193 714 193 1 co_n_6_M1
rlabel metal1 701 173 701 173 1 co_6_M1
rlabel metal1 612 186 612 186 1 zc1_n_5_M1
rlabel metal1 598 186 598 186 1 c1_5_M1
rlabel metal1 560 206 560 206 1 cn_5_M1
rlabel ntransistor 577 173 577 173 1 s_fa5_n_M1
rlabel metal1 488 211 488 211 1 bn_5_M1
rlabel ptransistor 484 195 484 195 1 an_5_M1
rlabel metal1 500 190 500 190 1 so_5_M1
rlabel metal1 387 190 387 190 1 co_5__M1
rlabel metal1 283 184 283 184 1 zc1_4_M1
rlabel metal1 269 184 269 184 1 c1_4_M1
rlabel ntransistor 248 171 248 171 1 s_fa4_n_M1
rlabel metal1 231 204 231 204 1 cn_1_M1
rlabel metal1 148 203 148 203 1 bn4_M1
rlabel ptransistor 155 193 155 193 1 an4_M1
rlabel metal1 171 188 171 188 1 so_4_M1
rlabel metal1 58 188 58 188 1 co_n4_M1
rlabel metal1 45 168 45 168 1 co_4_M1
rlabel metal1 154 118 154 118 1 a5_n_M1
rlabel metal1 491 124 491 124 1 c_fa5_M1
rlabel metal1 483 120 483 120 1 c_fa5_n_M1
rlabel metal1 810 123 810 123 1 c_fa6_n_M1
rlabel metal1 818 127 818 127 1 c_fa6_M1
rlabel metal1 511 30 511 30 1 q2b0_M1
rlabel metal1 520 29 520 29 1 q2b0_n_M1
rlabel m2contact 548 28 548 28 1 q2_M1
rlabel metal1 423 30 423 30 1 q2b1_M1
rlabel metal1 432 30 432 30 1 q2b1_n_M1
rlabel metal1 353 19 353 19 1 q2b2_n_M1
rlabel metal1 331 18 331 18 1 q2b2_M1
rlabel metal1 140 421 140 421 1 q0b2_n_M1
rlabel metal1 235 421 235 421 1 q0b1_M1
rlabel metal1 544 414 544 414 1 q1b0_n_M1
rlabel metal1 227 422 227 422 1 q0b1_n_M1
rlabel metal1 327 423 327 423 1 a0_M1
rlabel m2contact 1063 406 1063 406 1 en_bar_D1
rlabel metal1 1134 413 1134 413 1 D_bar_D1
rlabel metal1 1181 411 1181 411 1 out_n1_D1
rlabel ndiffusion 1162 394 1162 394 1 n1_D1
rlabel ndiffusion 1218 394 1218 394 1 n2_D1
rlabel metal1 1236 407 1236 407 1 out_n2_D1
rlabel ndiffusion 1274 394 1274 394 1 n3_D1
rlabel ndiffusion 1328 394 1328 394 1 n4_D1
rlabel m2contact 1345 410 1345 410 1 q_l1_bar_D1
rlabel m2contact 1349 353 1349 353 1 q_bar_D1
rlabel ndiffusion 1332 369 1332 369 1 n10_D1
rlabel metal1 1240 356 1240 356 1 out_n8_D1
rlabel ndiffusion 1222 369 1222 369 1 n8_D1
rlabel metal1 1185 352 1185 352 1 out_n7_D1
rlabel ndiffusion 1166 369 1166 369 1 n7_D1
rlabel polycontact 1156 349 1156 349 1 q_l1_D1
rlabel metal1 1138 353 1138 353 1 n6_D1
rlabel ndiffusion 1278 369 1278 369 1 n9_D1
rlabel m2contact 1295 345 1295 345 1 q_D1
rlabel m2contact 1345 265 1345 265 1 q_l1_bar_D2
rlabel metal1 1138 208 1138 208 1 n6_D2
rlabel polycontact 1156 204 1156 204 1 q_l1_D2
rlabel ndiffusion 1166 224 1166 224 1 n7_D2
rlabel metal1 1185 207 1185 207 1 out_n7__D2
rlabel ndiffusion 1222 224 1222 224 1 n8_D2
rlabel metal1 1240 211 1240 211 1 out_n8_D2
rlabel ndiffusion 1278 224 1278 224 1 n9_D2
rlabel m2contact 1295 200 1295 200 1 q_D2
rlabel ndiffusion 1332 224 1332 224 1 n10_D2
rlabel m2contact 1349 208 1349 208 1 q_bar_D2
rlabel ndiffusion 1328 249 1328 249 1 n4_D2
rlabel ndiffusion 1274 249 1274 249 1 n3_D2
rlabel metal1 1236 262 1236 262 1 out_n2_D2
rlabel ndiffusion 1218 249 1218 249 1 n2_D2
rlabel metal1 1181 266 1181 266 1 out_n1_D2
rlabel ndiffusion 1162 249 1162 249 1 n1_D2
rlabel metal1 1134 268 1134 268 1 D_bar_D2
rlabel m2contact 1063 261 1063 261 1 en_bar_D2
rlabel metal1 1137 66 1137 66 1 n6_D3
rlabel polycontact 1155 62 1155 62 1 q_l1_D3
rlabel ndiffusion 1165 82 1165 82 1 n7_D3
rlabel metal1 1184 65 1184 65 1 out_n7_D3
rlabel ndiffusion 1221 82 1221 82 1 n8_D3
rlabel m2contact 1294 58 1294 58 1 q_D3
rlabel metal1 1239 69 1239 69 1 out_n8_D3
rlabel ndiffusion 1277 82 1277 82 1 n9_D3
rlabel m2contact 1348 66 1348 66 1 q_bar_D3
rlabel m2contact 1344 123 1344 123 1 q_l1_bar_D3
rlabel ndiffusion 1327 107 1327 107 1 n4_D3
rlabel ndiffusion 1273 107 1273 107 1 n3_D3
rlabel metal1 1235 120 1235 120 1 out_n2_D3
rlabel ndiffusion 1217 107 1217 107 1 n2_D3
rlabel metal1 1180 124 1180 124 1 out_n1_D3
rlabel ndiffusion 1161 107 1161 107 1 n1_D3
rlabel metal1 1133 126 1133 126 1 D_bar_D3
rlabel m2contact 1062 119 1062 119 1 en_bar_D3
rlabel ndiffusion 1331 82 1331 82 1 n10
rlabel polycontact 1173 414 1173 414 1 en
rlabel polycontact 1381 269 1381 269 1 q_D1
rlabel polycontact 1394 270 1394 270 1 q_D1_n
rlabel polycontact 1382 209 1382 209 1 q_D2
rlabel polycontact 1395 209 1395 209 1 q_n_D2
rlabel polycontact 1382 130 1382 130 1 q_D3
rlabel polycontact 1394 130 1394 130 1 q_D3_n
rlabel metal2 1390 -459 1390 -459 7 q_D6
rlabel metal1 1160 -445 1160 -445 1 n6_D6
rlabel polycontact 1176 -449 1176 -449 1 q_l1_D6
rlabel metal1 1205 -446 1205 -446 1 out_n7_D6
rlabel ndiffusion 1186 -429 1186 -429 1 n7_D6
rlabel metal1 1260 -442 1260 -442 1 out_n8_D6
rlabel ndiffusion 1242 -429 1242 -429 1 n8_D6
rlabel m2contact 1315 -453 1315 -453 1 q_D6
rlabel ndiffusion 1298 -429 1298 -429 1 n9_D6
rlabel m2contact 1369 -445 1369 -445 1 q_bar_D6
rlabel ndiffusion 1352 -429 1352 -429 1 n10_D6
rlabel m2contact 1365 -388 1365 -388 1 q_l1_bar_D6
rlabel ndiffusion 1348 -404 1348 -404 1 n4_D6
rlabel ndiffusion 1294 -404 1294 -404 1 n3_D6
rlabel metal1 1256 -391 1256 -391 1 out_n2_D6
rlabel ndiffusion 1238 -404 1238 -404 1 n2_D6
rlabel ndiffusion 1182 -404 1182 -404 1 n1_D6
rlabel metal1 1201 -387 1201 -387 1 out_n1_D6
rlabel polycontact 1193 -384 1193 -384 1 en_D6
rlabel metal1 1154 -385 1154 -385 1 D_Bar_D6
rlabel m2contact 1083 -392 1083 -392 1 en_bar_D6
rlabel metal2 1388 -310 1388 -310 7 q_D5
rlabel metal1 1158 -303 1158 -303 1 n6_D5
rlabel polycontact 1175 -307 1175 -307 1 q_l1_D5
rlabel ndiffusion 1185 -287 1185 -287 1 n7_D5
rlabel metal1 1204 -304 1204 -304 1 out_n7_D5
rlabel ndiffusion 1241 -287 1241 -287 1 n8_D5
rlabel metal1 1259 -300 1259 -300 1 out_n8_D5
rlabel m2contact 1314 -311 1314 -311 1 q_D5
rlabel ndiffusion 1297 -287 1297 -287 1 n9_D5
rlabel metal1 1368 -295 1368 -295 1 q_bar_D5
rlabel ndiffusion 1351 -287 1351 -287 1 n10_D5
rlabel metal1 1364 -241 1364 -241 1 q_l1_bar_D5
rlabel ndiffusion 1347 -262 1347 -262 1 n4_D5
rlabel ndiffusion 1293 -262 1293 -262 1 n3_D5
rlabel metal1 1255 -249 1255 -249 1 out_n2_D5
rlabel ndiffusion 1237 -262 1237 -262 1 n2_D5
rlabel ndiffusion 1181 -262 1181 -262 1 n1_D5
rlabel metal1 1200 -245 1200 -245 1 out_n1_D5
rlabel polycontact 1192 -242 1192 -242 1 en_D5
rlabel metal1 1153 -243 1153 -243 1 D_bar_D5
rlabel m2contact 1082 -250 1082 -250 1 en_bar_D5
rlabel metal1 1202 -100 1202 -100 1 out_n1_D4
rlabel metal1 1159 -158 1159 -158 1 n6_D4
rlabel polycontact 1177 -162 1177 -162 1 q_l1_D4
rlabel ndiffusion 1187 -142 1187 -142 1 n7_D4
rlabel metal1 1206 -159 1206 -159 1 out_n7_D4
rlabel metal1 1261 -155 1261 -155 1 out_n8_D4
rlabel ndiffusion 1243 -142 1243 -142 1 n8_D4
rlabel ndiffusion 1299 -142 1299 -142 1 n9_D4
rlabel m2contact 1316 -166 1316 -166 1 q_D4
rlabel m2contact 1370 -158 1370 -158 1 q_bar_D4
rlabel ndiffusion 1353 -142 1353 -142 1 n10_D4
rlabel m2contact 1364 -102 1364 -102 1 q_l1_bar_D4
rlabel ndiffusion 1349 -117 1349 -117 1 n4_D4
rlabel ndiffusion 1295 -117 1295 -117 1 n3_D4
rlabel metal1 1257 -104 1257 -104 1 out_n2_D4
rlabel ndiffusion 1239 -117 1239 -117 1 n2_D4
rlabel ndiffusion 1183 -117 1183 -117 1 n1_D4
rlabel polycontact 1194 -97 1194 -97 1 en_D4
rlabel metal1 1155 -98 1155 -98 1 D_bar_D4
rlabel m2contact 1084 -105 1084 -105 1 en_bar_D4
rlabel m2contact 123 -81 123 -81 1 q0_M2
rlabel metal1 151 -85 151 -85 1 q0b2_n_M2
rlabel metal1 159 -89 159 -89 1 q0b2_M2
rlabel metal1 238 -84 238 -84 1 q0b1_n_M2
rlabel metal1 246 -85 246 -85 1 q0b1_M2
rlabel metal1 331 -82 331 -82 1 q0b0_n_M2
rlabel metal1 451 -76 451 -76 1 b2_M2
rlabel metal1 452 -116 452 -116 1 b0_M2
rlabel metal1 452 -97 452 -97 1 b1_M2
rlabel metal1 648 -71 648 -71 1 q1b1_M2
rlabel metal1 726 -82 726 -82 1 q1b2_M2
rlabel metal1 735 -82 735 -82 1 q1b2_n_M2
rlabel m2contact 762 -79 762 -79 1 q1_M2
rlabel metal1 951 -171 951 -171 1 zc1_n_3_M2
rlabel metal1 937 -171 937 -171 1 c1_3_M2
rlabel metal1 923 -167 923 -167 1 s_fa3_M2
rlabel ntransistor 916 -184 916 -184 1 s_fa3_n_M2
rlabel metal1 839 -167 839 -167 1 so_3_M2
rlabel metal1 726 -167 726 -167 1 co_n3_M2
rlabel metal1 713 -187 713 -187 1 co_3_M2
rlabel metal1 624 -174 624 -174 1 zc1_2_n_M2
rlabel metal1 610 -174 610 -174 1 c1_2_M2
rlabel pdcontact 586 -157 586 -157 1 s_fa2_M2
rlabel metal1 574 -174 574 -174 1 cn2_M2
rlabel ntransistor 589 -187 589 -187 1 son_2_M2
rlabel metal1 512 -170 512 -170 1 so_2_M2
rlabel polycontact 495 -173 495 -173 1 bn_2_M2
rlabel polycontact 504 -173 504 -173 1 an_2_M2
rlabel metal1 399 -171 399 -171 1 co_n2_M2
rlabel metal1 386 -190 386 -190 1 co_2_M2
rlabel metal1 295 -176 295 -176 1 zc1_n1_M2
rlabel metal1 281 -176 281 -176 1 c1_1_M2
rlabel ntransistor 260 -189 260 -189 1 a1_1_M2
rlabel metal1 183 -172 183 -172 1 so_1_M2
rlabel ntransistor 176 -188 176 -188 1 an_1_M2
rlabel metal1 171 -151 171 -151 1 bn_1_M1
rlabel metal1 57 -192 57 -192 1 co_1_M2
rlabel metal1 70 -172 70 -172 1 co_n1_M2
rlabel metal1 166 -244 166 -244 1 c_fa1_n_M2
rlabel metal1 174 -244 174 -244 1 c_fa1_M2
rlabel metal1 495 -240 495 -240 1 c_fa2_n_M2
rlabel metal1 503 -236 503 -236 1 c_fa2_M2
rlabel metal1 822 -237 822 -237 1 c_fa3_n_M2
rlabel metal1 830 -233 830 -233 1 c_fa3_M2
rlabel metal1 950 -317 950 -317 1 zc1_6_n_M2
rlabel metal1 936 -317 936 -317 1 c1_6_M2
rlabel ntransistor 915 -330 915 -330 1 s_fa_6_n_M2
rlabel metal1 898 -296 898 -296 1 cn_6_M2
rlabel metal1 838 -313 838 -313 1 so_6_M2
rlabel ptransistor 822 -308 822 -308 1 an_6_M2
rlabel metal1 783 -319 783 -319 1 bn_6_M2
rlabel metal1 725 -313 725 -313 1 co_n_6_M2
rlabel metal1 712 -333 712 -333 1 co_6_M2
rlabel ntransistor 588 -333 588 -333 1 s_fa_5_n_M2
rlabel metal1 499 -295 499 -295 1 bn_5_M2
rlabel ptransistor 495 -311 495 -311 1 an_5_M2
rlabel metal1 511 -316 511 -316 1 so_5_M2
rlabel metal1 294 -322 294 -322 1 zc1_4_M2
rlabel metal1 280 -322 280 -322 1 c1_4_M2
rlabel ntransistor 259 -335 259 -335 1 s_fa4_n_M2
rlabel metal1 242 -302 242 -302 1 cn_1_M2
rlabel metal1 159 -303 159 -303 1 bn4_M2
rlabel ptransistor 166 -313 166 -313 1 an4_M2
rlabel metal1 182 -318 182 -318 1 so_4_M2
rlabel metal1 69 -318 69 -318 1 co_n4_M2
rlabel metal1 56 -338 56 -338 1 co_4_M2
rlabel polycontact 165 -385 165 -385 1 a5_n_M2
rlabel metal1 494 -386 494 -386 1 c_fa5_n_M2
rlabel metal1 502 -382 502 -382 1 c_fa5_M2
rlabel metal1 821 -383 821 -383 1 c_fa6_n_M2
rlabel metal1 829 -379 829 -379 1 c_fa6_M2
rlabel metal1 364 -487 364 -487 1 q2b2_n_M2
rlabel metal1 342 -488 342 -488 1 q2b2_M2
rlabel metal1 434 -476 434 -476 1 q2b1_M2
rlabel metal1 443 -476 443 -476 1 q2b1_n_M2
rlabel m2contact 559 -478 559 -478 1 q2_M2
rlabel metal1 531 -477 531 -477 1 q2b0_n_M2
rlabel metal1 522 -476 522 -476 1 q2b0_M2
rlabel metal1 546 -78 546 -78 1 q1b0_M2
rlabel metal1 555 -92 555 -92 1 q1b0_n_M2
rlabel metal1 900 -149 900 -149 1 cn_3_M2
rlabel ptransistor 823 -162 823 -162 1 an3_M2
rlabel metal1 827 -146 827 -146 1 bn3_M2
rlabel metal1 398 -316 398 -316 1 co_5_M2
rlabel metal1 648 -93 648 -93 1 q1b1_n_M2
rlabel metal1 23 -86 23 -86 1 q0_M2
rlabel metal2 21 -38 21 -38 5 q1_M2
rlabel metal1 302 -478 303 -478 1 q2_M2
rlabel metal2 1388 -165 1388 -165 1 q_D4
rlabel metal1 1434 -268 1434 -268 1 buf_q_D4
rlabel polycontact 1426 -264 1426 -264 1 q_D4_n
rlabel polycontact 1428 -365 1429 -365 1 q_D5_n
rlabel metal1 1436 -361 1436 -361 1 buf_q_D5
rlabel polycontact 1430 -443 1430 -443 1 q_D6_n
rlabel metal1 1438 -446 1438 -446 1 buf_q_D6
rlabel metal1 1677 -487 1677 -487 7 n1_A1
rlabel metal1 1697 -500 1697 -500 7 n5_A1
rlabel metal1 1661 -430 1661 -430 7 b1_A1
rlabel metal1 1656 -386 1656 -386 7 bn_A1
rlabel metal1 1683 -429 1683 -429 7 b1n_A1
rlabel polycontact 1685 -414 1685 -414 7 a1_A1
rlabel metal1 1677 -374 1677 -374 7 xor1_A1
rlabel ndcontact 1693 -403 1693 -403 7 a1n_A1
rlabel metal1 1662 -314 1662 -314 7 n3_A1
rlabel metal1 1677 -290 1677 -290 7 s1_A1
rlabel metal1 1681 -276 1681 -276 7 c1_A1
rlabel metal1 1681 -262 1681 -262 7 zc1_n_A1
rlabel metal1 1685 -131 1685 -131 7 n9_n_A1
rlabel metal1 1705 -144 1705 -144 7 n9_A1
rlabel metal1 1668 -74 1668 -74 7 b2_A1
rlabel metal1 1691 -73 1691 -73 7 b2n_A1
rlabel metal1 1697 -66 1697 -66 7 a2_A1
rlabel ptransistor 1680 -34 1680 -34 7 a2n_A1
rlabel metal1 1685 -18 1685 -18 7 xor_2_A1
rlabel metal2 1665 2 1665 2 7 s2_A1
rlabel metal1 1668 43 1668 43 7 n6_A1
rlabel metal1 1685 66 1685 66 7 s3_A1
rlabel ntransistor 1702 59 1702 59 7 n7_A1
rlabel metal1 1689 80 1689 80 7 n8_A1
rlabel metal1 1689 94 1689 94 7 zc2_n_A1
rlabel metal1 1585 75 1585 75 7 n10_A1
rlabel metal1 1605 62 1605 62 7 n10_nA1
rlabel m2contact 1670 -193 1670 -193 7 s2_A1
rlabel ntransistor 1589 -44 1589 -44 7 a3n_A1
rlabel polycontact 1597 -11 1597 -11 7 a3_A1
rlabel metal1 1605 -51 1605 -51 7 xor_3_A1
rlabel polycontact 1602 -42 1602 -42 7 a3n_A1
rlabel metal1 1602 -27 1602 -27 7 b3n_A1
rlabel metal1 1621 5 1621 5 7 b3_A1
rlabel m2contact 1539 -42 1539 -42 7 c3_A1
rlabel metal1 1535 -34 1535 -34 7 cout3_n_A1
rlabel metal1 1755 -35 1755 -35 7 cout2_n_A1
rlabel metal1 1752 -27 1752 -27 7 c2_A1
rlabel ntransistor 1588 -128 1588 -128 7 n11_A1
rlabel metal1 1605 -135 1605 -135 7 s4_a1
rlabel metal1 1621 -107 1621 -107 7 n12_A1
rlabel metal2 1625 -87 1625 -87 7 c2_A1
rlabel metal1 1601 -149 1601 -149 7 n13_A1
rlabel metal1 1601 -163 1601 -163 7 zc3_n_A1
rlabel metal1 1747 -391 1747 -391 7 cout_n_A1
rlabel metal1 1743 -383 1743 -383 7 s2_A1
rlabel metal1 1726 -503 1726 -503 7 co_A1
rlabel metal1 1729 -472 1729 -472 7 n2_A1
rlabel polycontact 1735 -439 1735 -439 7 son_A1
rlabel polycontact 1745 -445 1745 -445 7 con_A1
rlabel metal1 1742 -431 1742 -431 7 so_A1
rlabel metal1 1746 -463 1746 -463 7 b_A1
rlabel polycontact 1742 -487 1742 -487 7 a_A1
rlabel metal1 1599 197 1599 197 7 zc5_n_A1
rlabel metal1 1599 211 1599 211 7 n21_A1
rlabel ntransistor 1586 232 1586 232 7 n19_A1
rlabel metal1 1603 225 1603 225 7 s6_A1
rlabel metal1 1619 253 1619 253 7 n20_A1
rlabel metal2 1623 273 1623 273 7 c4_A1
rlabel ntransistor 1587 316 1587 316 7 a5n_A1
rlabel polycontact 1595 349 1595 349 7 a5_A1
rlabel metal1 1603 309 1603 309 7 xor_5_A1
rlabel metal1 1600 333 1600 333 7 b5n_A1
rlabel metal1 1619 365 1619 365 7 b5_A1
rlabel metal1 1583 435 1583 435 7 n18_A1
rlabel metal2 1668 167 1668 167 7 c3_A1
rlabel metal1 1683 229 1683 229 7 n17n_A1
rlabel metal1 1703 216 1703 216 7 n17_A1
rlabel metal1 1666 286 1666 286 7 b4_A1
rlabel metal1 1689 287 1689 287 7 b4n_A1
rlabel metal1 1695 294 1695 294 7 a4_A1
rlabel ptransistor 1678 326 1678 326 7 a4n_A1
rlabel metal1 1683 342 1683 342 7 xor_4_A1
rlabel metal2 1663 362 1663 362 7 c3_A1
rlabel metal1 1666 403 1666 403 7 n14_A1
rlabel metal1 1683 426 1683 426 7 s5_A1
rlabel ntransistor 1700 419 1700 419 7 n15_A1
rlabel metal1 1687 440 1687 440 7 n16_A1
rlabel metal1 1687 454 1687 454 7 zc4_n_A1
rlabel metal1 1749 333 1749 333 7 c4_A1
rlabel metal1 1753 325 1753 325 7 cout4n_A1
rlabel metal1 1537 318 1537 318 7 c5_A1
rlabel metal1 1533 326 1533 326 7 cout5_n_A1
rlabel metal1 1603 422 1603 422 7 n18_nA1
rlabel metal2 1677 -557 1677 -557 7 a1_A1
rlabel metal2 1799 -561 1799 -561 7 b2_A1
rlabel metal1 1548 -252 1548 -252 7 a3_A1
rlabel metal1 1558 -253 1558 -253 7 b3_A1
rlabel metal2 1810 -560 1810 -560 7 a4_A1
rlabel metal2 1825 -563 1825 -563 7 b4_A1
rlabel metal2 1508 -144 1508 -144 7 b5_A1
rlabel metal2 1491 -149 1491 -149 3 a5_A1
rlabel polycontact 1680 -298 1680 -298 7 n4_A1
rlabel metal2 1491 482 1491 482 4 s1_A1
rlabel metal1 1832 491 1832 491 7 so_A1
rlabel metal2 1797 498 1797 498 5 s3_A1
rlabel metal1 1817 497 1817 497 7 s1_A1
rlabel metal2 1783 500 1783 500 5 s5_A1
rlabel metal2 1773 500 1773 500 5 s6_A1
rlabel metal2 1509 491 1509 491 7 c5_A1
rlabel metal2 1560 492 1560 492 7 s4_A1
rlabel metal2 1767 -560 1767 -560 1 a_A1
rlabel polysilicon 1772 -561 1772 -561 1 b_A1
rlabel metal2 1786 -559 1786 -559 1 a2_A1
rlabel polycontact 904 336 904 336 1 s_fa3_n_M1
rlabel polycontact 154 331 154 331 1 bn_n_M1
rlabel metal1 571 -300 571 -300 1 cn_5_M2
rlabel metal1 609 -320 609 -320 1 c1_5_M2
rlabel metal1 623 -320 623 -320 1 zc1_n_5_M2
rlabel metal1 206 446 206 446 1 vss
rlabel metal1 140 368 140 368 1 vdd
rlabel metal2 1664 -558 1664 -558 1 b1_A1
<< end >>
