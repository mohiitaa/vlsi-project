magic
tech scmos
timestamp 1523040320
<< pwell >>
rect 110 457 128 461
rect 108 453 128 457
rect 108 417 156 453
rect 195 417 243 453
rect 288 417 336 453
rect 528 419 576 455
rect 621 419 669 455
rect 708 419 756 455
rect 37 294 180 330
rect 192 294 310 330
rect 366 296 509 332
rect 521 296 639 332
rect 693 299 836 335
rect 848 299 966 335
rect 123 268 171 294
rect 452 270 500 296
rect 779 273 827 299
rect 36 148 179 184
rect 191 148 309 184
rect 365 150 508 186
rect 520 150 638 186
rect 692 153 835 189
rect 847 153 965 189
rect 122 122 170 148
rect 451 124 499 150
rect 778 127 826 153
rect 323 0 371 36
rect 416 0 464 36
rect 503 0 551 36
<< nwell >>
rect 108 374 156 417
rect 195 374 243 417
rect 288 374 336 417
rect 528 382 576 419
rect 621 382 669 419
rect 528 379 669 382
rect 524 376 669 379
rect 1005 421 1184 447
rect 1197 421 1238 447
rect 1253 421 1294 447
rect 1307 421 1348 447
rect 708 388 756 419
rect 708 379 769 388
rect 708 376 836 379
rect 37 330 180 374
rect 192 373 336 374
rect 192 330 310 373
rect 366 332 509 376
rect 521 362 836 376
rect 521 332 639 362
rect 693 335 836 362
rect 848 335 966 379
rect 1101 316 1188 342
rect 1201 316 1242 342
rect 1257 316 1298 342
rect 1311 316 1352 342
rect 123 261 171 268
rect 452 263 500 270
rect 1005 276 1184 302
rect 1197 276 1238 302
rect 1253 276 1294 302
rect 1307 276 1348 302
rect 779 266 827 273
rect 119 248 171 261
rect 448 250 500 263
rect 775 253 827 266
rect 123 232 171 248
rect 452 234 500 250
rect 779 240 827 253
rect 112 228 178 232
rect 442 230 508 234
rect 750 233 861 240
rect 36 184 179 228
rect 191 184 309 228
rect 365 186 508 230
rect 520 186 638 230
rect 692 224 965 233
rect 692 189 835 224
rect 847 189 965 224
rect 1101 171 1188 197
rect 1201 171 1242 197
rect 1257 171 1298 197
rect 1311 171 1352 197
rect 1040 160 1059 162
rect 122 115 170 122
rect 451 117 499 124
rect 1004 134 1183 160
rect 1196 134 1237 160
rect 1252 134 1293 160
rect 1306 134 1347 160
rect 778 120 826 127
rect 118 102 170 115
rect 447 104 499 117
rect 774 107 826 120
rect 122 78 170 102
rect 451 94 499 104
rect 325 80 557 94
rect 778 83 826 107
rect 323 77 557 80
rect 323 36 371 77
rect 416 36 464 77
rect 503 36 551 77
rect 1100 29 1187 55
rect 1200 29 1241 55
rect 1256 29 1297 55
rect 1310 29 1351 55
<< polysilicon >>
rect 121 436 123 441
rect 128 436 130 441
rect 141 434 143 438
rect 208 436 210 441
rect 215 436 217 441
rect 228 434 230 438
rect 301 436 303 441
rect 308 436 310 441
rect 321 434 323 438
rect 541 436 543 440
rect 554 438 556 443
rect 561 438 563 443
rect 634 436 636 440
rect 647 438 649 443
rect 654 438 656 443
rect 721 436 723 440
rect 734 438 736 443
rect 741 438 743 443
rect 1042 434 1044 436
rect 1114 434 1116 440
rect 1153 434 1155 440
rect 1174 434 1176 440
rect 1207 434 1209 440
rect 1228 434 1230 440
rect 1263 434 1265 440
rect 1284 434 1286 440
rect 1317 434 1319 440
rect 1338 434 1340 440
rect 121 412 123 425
rect 128 420 130 425
rect 141 420 143 425
rect 127 419 133 420
rect 127 415 128 419
rect 132 415 133 419
rect 127 414 133 415
rect 137 419 143 420
rect 137 415 138 419
rect 142 415 143 419
rect 137 414 143 415
rect 117 411 123 412
rect 117 407 118 411
rect 122 407 123 411
rect 117 406 123 407
rect 121 403 123 406
rect 131 403 133 414
rect 141 410 143 414
rect 208 412 210 425
rect 215 420 217 425
rect 228 420 230 425
rect 214 419 220 420
rect 214 415 215 419
rect 219 415 220 419
rect 214 414 220 415
rect 224 419 230 420
rect 224 415 225 419
rect 229 415 230 419
rect 224 414 230 415
rect 204 411 210 412
rect 204 407 205 411
rect 209 407 210 411
rect 204 406 210 407
rect 208 403 210 406
rect 218 403 220 414
rect 228 410 230 414
rect 301 412 303 425
rect 308 420 310 425
rect 321 420 323 425
rect 307 419 313 420
rect 307 415 308 419
rect 312 415 313 419
rect 307 414 313 415
rect 317 419 323 420
rect 317 415 318 419
rect 322 415 323 419
rect 317 414 323 415
rect 297 411 303 412
rect 121 385 123 390
rect 131 385 133 390
rect 141 388 143 392
rect 297 407 298 411
rect 302 407 303 411
rect 297 406 303 407
rect 301 403 303 406
rect 311 403 313 414
rect 321 410 323 414
rect 541 422 543 427
rect 554 422 556 427
rect 541 421 547 422
rect 541 417 542 421
rect 546 417 547 421
rect 541 416 547 417
rect 551 421 557 422
rect 551 417 552 421
rect 556 417 557 421
rect 551 416 557 417
rect 541 412 543 416
rect 208 385 210 390
rect 218 385 220 390
rect 228 388 230 392
rect 551 405 553 416
rect 561 414 563 427
rect 634 422 636 427
rect 647 422 649 427
rect 634 421 640 422
rect 634 417 635 421
rect 639 417 640 421
rect 634 416 640 417
rect 644 421 650 422
rect 644 417 645 421
rect 649 417 650 421
rect 644 416 650 417
rect 561 413 567 414
rect 561 409 562 413
rect 566 409 567 413
rect 634 412 636 416
rect 561 408 567 409
rect 561 405 563 408
rect 301 385 303 390
rect 311 385 313 390
rect 321 388 323 392
rect 541 390 543 394
rect 644 405 646 416
rect 654 414 656 427
rect 721 422 723 427
rect 734 422 736 427
rect 721 421 727 422
rect 721 417 722 421
rect 726 417 727 421
rect 721 416 727 417
rect 731 421 737 422
rect 731 417 732 421
rect 736 417 737 421
rect 731 416 737 417
rect 654 413 660 414
rect 654 409 655 413
rect 659 409 660 413
rect 721 412 723 416
rect 654 408 660 409
rect 654 405 656 408
rect 551 387 553 392
rect 561 387 563 392
rect 634 390 636 394
rect 731 405 733 416
rect 741 414 743 427
rect 1042 417 1044 428
rect 741 413 747 414
rect 1114 416 1116 428
rect 1153 416 1155 428
rect 1174 416 1176 428
rect 1207 416 1209 428
rect 1228 416 1230 428
rect 1263 416 1265 428
rect 1284 416 1286 428
rect 1317 416 1319 428
rect 1338 416 1340 428
rect 741 409 742 413
rect 746 409 747 413
rect 741 408 747 409
rect 741 405 743 408
rect 644 387 646 392
rect 654 387 656 392
rect 721 390 723 394
rect 1042 395 1044 413
rect 1154 412 1155 416
rect 1175 412 1176 416
rect 1208 412 1209 416
rect 1229 412 1230 416
rect 1264 412 1265 416
rect 1285 412 1286 416
rect 1318 412 1319 416
rect 1339 412 1340 416
rect 731 387 733 392
rect 741 387 743 392
rect 1042 389 1044 392
rect 1114 394 1116 412
rect 1153 397 1155 412
rect 1174 397 1176 412
rect 1207 397 1209 412
rect 1228 397 1230 412
rect 1263 397 1265 412
rect 1284 397 1286 412
rect 1317 397 1319 412
rect 1338 397 1340 412
rect 1114 388 1116 391
rect 1153 388 1155 391
rect 1174 388 1176 391
rect 1207 388 1209 391
rect 1228 388 1230 391
rect 1263 388 1265 391
rect 1284 388 1286 391
rect 1317 388 1319 391
rect 1338 388 1340 391
rect 129 364 131 368
rect 53 356 59 357
rect 43 348 45 353
rect 53 352 54 356
rect 58 352 59 356
rect 53 351 59 352
rect 53 346 55 351
rect 63 346 65 351
rect 114 348 120 349
rect 114 344 115 348
rect 119 344 120 348
rect 114 343 120 344
rect 43 333 45 336
rect 53 333 55 336
rect 43 332 49 333
rect 43 328 44 332
rect 48 328 49 332
rect 53 330 57 333
rect 43 327 49 328
rect 43 319 45 327
rect 55 316 57 330
rect 63 325 65 336
rect 118 334 120 343
rect 165 364 167 368
rect 213 364 215 368
rect 145 355 147 359
rect 155 355 157 359
rect 198 348 204 349
rect 198 344 199 348
rect 203 344 204 348
rect 198 343 204 344
rect 129 334 131 337
rect 145 334 147 337
rect 155 334 157 337
rect 165 334 167 337
rect 118 332 131 334
rect 137 332 147 334
rect 151 333 157 334
rect 62 324 68 325
rect 121 324 123 332
rect 137 328 139 332
rect 151 329 152 333
rect 156 329 157 333
rect 151 328 157 329
rect 161 333 167 334
rect 161 329 162 333
rect 166 329 167 333
rect 202 334 204 343
rect 249 364 251 368
rect 229 355 231 359
rect 239 355 241 359
rect 458 366 460 370
rect 382 358 388 359
rect 285 356 291 357
rect 275 348 277 353
rect 285 352 286 356
rect 290 352 291 356
rect 285 351 291 352
rect 213 334 215 337
rect 229 334 231 337
rect 239 334 241 337
rect 249 334 251 337
rect 285 346 287 351
rect 295 346 297 351
rect 372 350 374 355
rect 382 354 383 358
rect 387 354 388 358
rect 382 353 388 354
rect 382 348 384 353
rect 392 348 394 353
rect 443 350 449 351
rect 443 346 444 350
rect 448 346 449 350
rect 443 345 449 346
rect 202 332 215 334
rect 221 332 231 334
rect 235 333 241 334
rect 161 328 167 329
rect 130 327 139 328
rect 62 320 63 324
rect 67 320 68 324
rect 62 319 68 320
rect 62 316 64 319
rect 43 309 45 313
rect 130 323 131 327
rect 135 323 139 327
rect 155 324 157 328
rect 130 322 139 323
rect 137 319 139 322
rect 147 319 149 324
rect 155 322 159 324
rect 157 319 159 322
rect 164 319 166 328
rect 205 324 207 332
rect 221 328 223 332
rect 235 329 236 333
rect 240 329 241 333
rect 235 328 241 329
rect 245 333 251 334
rect 245 329 246 333
rect 250 329 251 333
rect 245 328 251 329
rect 275 333 277 336
rect 285 333 287 336
rect 275 332 281 333
rect 275 328 276 332
rect 280 328 281 332
rect 285 330 289 333
rect 214 327 223 328
rect 121 312 123 315
rect 121 310 126 312
rect 55 302 57 307
rect 62 302 64 307
rect 124 302 126 310
rect 137 306 139 310
rect 147 302 149 310
rect 214 323 215 327
rect 219 323 223 327
rect 239 324 241 328
rect 214 322 223 323
rect 221 319 223 322
rect 231 319 233 324
rect 239 322 243 324
rect 241 319 243 322
rect 248 319 250 328
rect 275 327 281 328
rect 275 319 277 327
rect 205 312 207 315
rect 205 310 210 312
rect 157 302 159 307
rect 164 302 166 307
rect 124 300 149 302
rect 208 302 210 310
rect 221 306 223 310
rect 231 302 233 310
rect 287 316 289 330
rect 295 325 297 336
rect 372 335 374 338
rect 382 335 384 338
rect 372 334 378 335
rect 372 330 373 334
rect 377 330 378 334
rect 382 332 386 335
rect 372 329 378 330
rect 294 324 300 325
rect 294 320 295 324
rect 299 320 300 324
rect 372 321 374 329
rect 294 319 300 320
rect 294 316 296 319
rect 275 309 277 313
rect 384 318 386 332
rect 392 327 394 338
rect 447 336 449 345
rect 494 366 496 370
rect 542 366 544 370
rect 474 357 476 361
rect 484 357 486 361
rect 527 350 533 351
rect 527 346 528 350
rect 532 346 533 350
rect 527 345 533 346
rect 458 336 460 339
rect 474 336 476 339
rect 484 336 486 339
rect 494 336 496 339
rect 447 334 460 336
rect 466 334 476 336
rect 480 335 486 336
rect 391 326 397 327
rect 450 326 452 334
rect 466 330 468 334
rect 480 331 481 335
rect 485 331 486 335
rect 480 330 486 331
rect 490 335 496 336
rect 490 331 491 335
rect 495 331 496 335
rect 531 336 533 345
rect 578 366 580 370
rect 558 357 560 361
rect 568 357 570 361
rect 785 369 787 373
rect 709 361 715 362
rect 614 358 620 359
rect 604 350 606 355
rect 614 354 615 358
rect 619 354 620 358
rect 614 353 620 354
rect 699 353 701 358
rect 709 357 710 361
rect 714 357 715 361
rect 709 356 715 357
rect 542 336 544 339
rect 558 336 560 339
rect 568 336 570 339
rect 578 336 580 339
rect 614 348 616 353
rect 624 348 626 353
rect 709 351 711 356
rect 719 351 721 356
rect 770 353 776 354
rect 770 349 771 353
rect 775 349 776 353
rect 770 348 776 349
rect 699 338 701 341
rect 709 338 711 341
rect 531 334 544 336
rect 550 334 560 336
rect 564 335 570 336
rect 490 330 496 331
rect 459 329 468 330
rect 391 322 392 326
rect 396 322 397 326
rect 391 321 397 322
rect 391 318 393 321
rect 372 311 374 315
rect 459 325 460 329
rect 464 325 468 329
rect 484 326 486 330
rect 459 324 468 325
rect 466 321 468 324
rect 476 321 478 326
rect 484 324 488 326
rect 486 321 488 324
rect 493 321 495 330
rect 534 326 536 334
rect 550 330 552 334
rect 564 331 565 335
rect 569 331 570 335
rect 564 330 570 331
rect 574 335 580 336
rect 574 331 575 335
rect 579 331 580 335
rect 574 330 580 331
rect 604 335 606 338
rect 614 335 616 338
rect 604 334 610 335
rect 604 330 605 334
rect 609 330 610 334
rect 614 332 618 335
rect 543 329 552 330
rect 450 314 452 317
rect 450 312 455 314
rect 241 302 243 307
rect 248 302 250 307
rect 208 300 233 302
rect 287 302 289 307
rect 294 302 296 307
rect 384 304 386 309
rect 391 304 393 309
rect 453 304 455 312
rect 466 308 468 312
rect 476 304 478 312
rect 543 325 544 329
rect 548 325 552 329
rect 568 326 570 330
rect 543 324 552 325
rect 550 321 552 324
rect 560 321 562 326
rect 568 324 572 326
rect 570 321 572 324
rect 577 321 579 330
rect 604 329 610 330
rect 604 321 606 329
rect 534 314 536 317
rect 534 312 539 314
rect 486 304 488 309
rect 493 304 495 309
rect 453 302 478 304
rect 537 304 539 312
rect 550 308 552 312
rect 560 304 562 312
rect 616 318 618 332
rect 624 327 626 338
rect 699 337 705 338
rect 699 333 700 337
rect 704 333 705 337
rect 709 335 713 338
rect 699 332 705 333
rect 623 326 629 327
rect 623 322 624 326
rect 628 322 629 326
rect 699 324 701 332
rect 623 321 629 322
rect 623 318 625 321
rect 711 321 713 335
rect 719 330 721 341
rect 774 339 776 348
rect 821 369 823 373
rect 869 369 871 373
rect 801 360 803 364
rect 811 360 813 364
rect 854 353 860 354
rect 854 349 855 353
rect 859 349 860 353
rect 854 348 860 349
rect 785 339 787 342
rect 801 339 803 342
rect 811 339 813 342
rect 821 339 823 342
rect 774 337 787 339
rect 793 337 803 339
rect 807 338 813 339
rect 718 329 724 330
rect 777 329 779 337
rect 793 333 795 337
rect 807 334 808 338
rect 812 334 813 338
rect 807 333 813 334
rect 817 338 823 339
rect 817 334 818 338
rect 822 334 823 338
rect 858 339 860 348
rect 905 369 907 373
rect 1118 372 1120 375
rect 1157 372 1159 375
rect 1178 372 1180 375
rect 1211 372 1213 375
rect 1232 372 1234 375
rect 1267 372 1269 375
rect 1288 372 1290 375
rect 1321 372 1323 375
rect 1342 372 1344 375
rect 885 360 887 364
rect 895 360 897 364
rect 941 361 947 362
rect 931 353 933 358
rect 941 357 942 361
rect 946 357 947 361
rect 941 356 947 357
rect 869 339 871 342
rect 885 339 887 342
rect 895 339 897 342
rect 905 339 907 342
rect 941 351 943 356
rect 951 351 953 356
rect 1118 351 1120 369
rect 1157 351 1159 366
rect 1178 351 1180 366
rect 1211 351 1213 366
rect 1232 351 1234 366
rect 1267 351 1269 366
rect 1288 351 1290 366
rect 1321 351 1323 366
rect 1342 351 1344 366
rect 1158 347 1159 351
rect 1179 347 1180 351
rect 1212 347 1213 351
rect 1233 347 1234 351
rect 1268 347 1269 351
rect 1289 347 1290 351
rect 1322 347 1323 351
rect 1343 347 1344 351
rect 858 337 871 339
rect 877 337 887 339
rect 891 338 897 339
rect 817 333 823 334
rect 786 332 795 333
rect 718 325 719 329
rect 723 325 724 329
rect 718 324 724 325
rect 718 321 720 324
rect 604 311 606 315
rect 699 314 701 318
rect 786 328 787 332
rect 791 328 795 332
rect 811 329 813 333
rect 786 327 795 328
rect 793 324 795 327
rect 803 324 805 329
rect 811 327 815 329
rect 813 324 815 327
rect 820 324 822 333
rect 861 329 863 337
rect 877 333 879 337
rect 891 334 892 338
rect 896 334 897 338
rect 891 333 897 334
rect 901 338 907 339
rect 901 334 902 338
rect 906 334 907 338
rect 901 333 907 334
rect 931 338 933 341
rect 941 338 943 341
rect 931 337 937 338
rect 931 333 932 337
rect 936 333 937 337
rect 941 335 945 338
rect 870 332 879 333
rect 777 317 779 320
rect 777 315 782 317
rect 570 304 572 309
rect 577 304 579 309
rect 537 302 562 304
rect 616 304 618 309
rect 623 304 625 309
rect 711 307 713 312
rect 718 307 720 312
rect 780 307 782 315
rect 793 311 795 315
rect 803 307 805 315
rect 870 328 871 332
rect 875 328 879 332
rect 895 329 897 333
rect 870 327 879 328
rect 877 324 879 327
rect 887 324 889 329
rect 895 327 899 329
rect 897 324 899 327
rect 904 324 906 333
rect 931 332 937 333
rect 931 324 933 332
rect 861 317 863 320
rect 861 315 866 317
rect 813 307 815 312
rect 820 307 822 312
rect 780 305 805 307
rect 864 307 866 315
rect 877 311 879 315
rect 887 307 889 315
rect 943 321 945 335
rect 951 330 953 341
rect 1118 335 1120 347
rect 1157 335 1159 347
rect 1178 335 1180 347
rect 1211 335 1213 347
rect 1232 335 1234 347
rect 1267 335 1269 347
rect 1288 335 1290 347
rect 1321 335 1323 347
rect 1342 335 1344 347
rect 950 329 956 330
rect 950 325 951 329
rect 955 325 956 329
rect 950 324 956 325
rect 950 321 952 324
rect 1118 323 1120 329
rect 1157 323 1159 329
rect 1178 323 1180 329
rect 1211 323 1213 329
rect 1232 323 1234 329
rect 1267 323 1269 329
rect 1288 323 1290 329
rect 1321 323 1323 329
rect 1342 323 1344 329
rect 931 314 933 318
rect 897 307 899 312
rect 904 307 906 312
rect 864 305 889 307
rect 943 307 945 312
rect 950 307 952 312
rect 136 285 138 289
rect 146 285 148 289
rect 156 285 158 289
rect 465 287 467 291
rect 475 287 477 291
rect 485 287 487 291
rect 792 290 794 294
rect 802 290 804 294
rect 812 290 814 294
rect 1042 289 1044 291
rect 136 271 138 279
rect 132 270 138 271
rect 146 270 148 279
rect 156 270 158 279
rect 465 273 467 281
rect 132 266 133 270
rect 137 266 138 270
rect 152 269 158 270
rect 132 265 138 266
rect 136 252 138 265
rect 146 263 148 266
rect 152 265 153 269
rect 157 265 158 269
rect 461 272 467 273
rect 475 272 477 281
rect 485 272 487 281
rect 792 276 794 284
rect 461 268 462 272
rect 466 268 467 272
rect 481 271 487 272
rect 461 267 467 268
rect 152 264 158 265
rect 142 262 148 263
rect 142 258 143 262
rect 147 258 148 262
rect 142 257 148 258
rect 143 252 145 257
rect 156 255 158 264
rect 465 254 467 267
rect 475 265 477 268
rect 481 267 482 271
rect 486 267 487 271
rect 788 275 794 276
rect 802 275 804 284
rect 812 275 814 284
rect 1114 289 1116 295
rect 1153 289 1155 295
rect 1174 289 1176 295
rect 1207 289 1209 295
rect 1228 289 1230 295
rect 1263 289 1265 295
rect 1284 289 1286 295
rect 1317 289 1319 295
rect 1338 289 1340 295
rect 788 271 789 275
rect 793 271 794 275
rect 808 274 814 275
rect 788 270 794 271
rect 481 266 487 267
rect 471 264 477 265
rect 471 260 472 264
rect 476 260 477 264
rect 471 259 477 260
rect 472 254 474 259
rect 485 257 487 266
rect 792 257 794 270
rect 802 268 804 271
rect 808 270 809 274
rect 813 270 814 274
rect 1042 272 1044 283
rect 808 269 814 270
rect 798 267 804 268
rect 798 263 799 267
rect 803 263 804 267
rect 798 262 804 263
rect 799 257 801 262
rect 812 260 814 269
rect 1114 271 1116 283
rect 1153 271 1155 283
rect 1174 271 1176 283
rect 1207 271 1209 283
rect 1228 271 1230 283
rect 1263 271 1265 283
rect 1284 271 1286 283
rect 1317 271 1319 283
rect 1338 271 1340 283
rect 156 239 158 243
rect 485 241 487 245
rect 812 244 814 248
rect 1042 250 1044 268
rect 1154 267 1155 271
rect 1175 267 1176 271
rect 1208 267 1209 271
rect 1229 267 1230 271
rect 1264 267 1265 271
rect 1285 267 1286 271
rect 1318 267 1319 271
rect 1339 267 1340 271
rect 1042 244 1044 247
rect 1114 249 1116 267
rect 1153 252 1155 267
rect 1174 252 1176 267
rect 1207 252 1209 267
rect 1228 252 1230 267
rect 1263 252 1265 267
rect 1284 252 1286 267
rect 1317 252 1319 267
rect 1338 252 1340 267
rect 1114 243 1116 246
rect 1153 243 1155 246
rect 1174 243 1176 246
rect 1207 243 1209 246
rect 1228 243 1230 246
rect 1263 243 1265 246
rect 1284 243 1286 246
rect 1317 243 1319 246
rect 1338 243 1340 246
rect 136 230 138 234
rect 143 230 145 234
rect 465 232 467 236
rect 472 232 474 236
rect 792 235 794 239
rect 799 235 801 239
rect 1118 227 1120 230
rect 1157 227 1159 230
rect 1178 227 1180 230
rect 1211 227 1213 230
rect 1232 227 1234 230
rect 1267 227 1269 230
rect 1288 227 1290 230
rect 1321 227 1323 230
rect 1342 227 1344 230
rect 128 218 130 222
rect 52 210 58 211
rect 42 202 44 207
rect 52 206 53 210
rect 57 206 58 210
rect 52 205 58 206
rect 52 200 54 205
rect 62 200 64 205
rect 113 202 119 203
rect 113 198 114 202
rect 118 198 119 202
rect 113 197 119 198
rect 42 187 44 190
rect 52 187 54 190
rect 42 186 48 187
rect 42 182 43 186
rect 47 182 48 186
rect 52 184 56 187
rect 42 181 48 182
rect 42 173 44 181
rect 54 170 56 184
rect 62 179 64 190
rect 117 188 119 197
rect 164 218 166 222
rect 212 218 214 222
rect 144 209 146 213
rect 154 209 156 213
rect 197 202 203 203
rect 197 198 198 202
rect 202 198 203 202
rect 197 197 203 198
rect 128 188 130 191
rect 144 188 146 191
rect 154 188 156 191
rect 164 188 166 191
rect 117 186 130 188
rect 136 186 146 188
rect 150 187 156 188
rect 61 178 67 179
rect 120 178 122 186
rect 136 182 138 186
rect 150 183 151 187
rect 155 183 156 187
rect 150 182 156 183
rect 160 187 166 188
rect 160 183 161 187
rect 165 183 166 187
rect 201 188 203 197
rect 248 218 250 222
rect 228 209 230 213
rect 238 209 240 213
rect 457 220 459 224
rect 381 212 387 213
rect 284 210 290 211
rect 274 202 276 207
rect 284 206 285 210
rect 289 206 290 210
rect 284 205 290 206
rect 212 188 214 191
rect 228 188 230 191
rect 238 188 240 191
rect 248 188 250 191
rect 284 200 286 205
rect 294 200 296 205
rect 371 204 373 209
rect 381 208 382 212
rect 386 208 387 212
rect 381 207 387 208
rect 381 202 383 207
rect 391 202 393 207
rect 442 204 448 205
rect 442 200 443 204
rect 447 200 448 204
rect 442 199 448 200
rect 201 186 214 188
rect 220 186 230 188
rect 234 187 240 188
rect 160 182 166 183
rect 129 181 138 182
rect 61 174 62 178
rect 66 174 67 178
rect 61 173 67 174
rect 61 170 63 173
rect 42 163 44 167
rect 129 177 130 181
rect 134 177 138 181
rect 154 178 156 182
rect 129 176 138 177
rect 136 173 138 176
rect 146 173 148 178
rect 154 176 158 178
rect 156 173 158 176
rect 163 173 165 182
rect 204 178 206 186
rect 220 182 222 186
rect 234 183 235 187
rect 239 183 240 187
rect 234 182 240 183
rect 244 187 250 188
rect 244 183 245 187
rect 249 183 250 187
rect 244 182 250 183
rect 274 187 276 190
rect 284 187 286 190
rect 274 186 280 187
rect 274 182 275 186
rect 279 182 280 186
rect 284 184 288 187
rect 213 181 222 182
rect 120 166 122 169
rect 120 164 125 166
rect 54 156 56 161
rect 61 156 63 161
rect 123 156 125 164
rect 136 160 138 164
rect 146 156 148 164
rect 213 177 214 181
rect 218 177 222 181
rect 238 178 240 182
rect 213 176 222 177
rect 220 173 222 176
rect 230 173 232 178
rect 238 176 242 178
rect 240 173 242 176
rect 247 173 249 182
rect 274 181 280 182
rect 274 173 276 181
rect 204 166 206 169
rect 204 164 209 166
rect 156 156 158 161
rect 163 156 165 161
rect 123 154 148 156
rect 207 156 209 164
rect 220 160 222 164
rect 230 156 232 164
rect 286 170 288 184
rect 294 179 296 190
rect 371 189 373 192
rect 381 189 383 192
rect 371 188 377 189
rect 371 184 372 188
rect 376 184 377 188
rect 381 186 385 189
rect 371 183 377 184
rect 293 178 299 179
rect 293 174 294 178
rect 298 174 299 178
rect 371 175 373 183
rect 293 173 299 174
rect 293 170 295 173
rect 274 163 276 167
rect 383 172 385 186
rect 391 181 393 192
rect 446 190 448 199
rect 493 220 495 224
rect 541 220 543 224
rect 473 211 475 215
rect 483 211 485 215
rect 526 204 532 205
rect 526 200 527 204
rect 531 200 532 204
rect 526 199 532 200
rect 457 190 459 193
rect 473 190 475 193
rect 483 190 485 193
rect 493 190 495 193
rect 446 188 459 190
rect 465 188 475 190
rect 479 189 485 190
rect 390 180 396 181
rect 449 180 451 188
rect 465 184 467 188
rect 479 185 480 189
rect 484 185 485 189
rect 479 184 485 185
rect 489 189 495 190
rect 489 185 490 189
rect 494 185 495 189
rect 530 190 532 199
rect 577 220 579 224
rect 557 211 559 215
rect 567 211 569 215
rect 784 223 786 227
rect 708 215 714 216
rect 613 212 619 213
rect 603 204 605 209
rect 613 208 614 212
rect 618 208 619 212
rect 613 207 619 208
rect 698 207 700 212
rect 708 211 709 215
rect 713 211 714 215
rect 708 210 714 211
rect 541 190 543 193
rect 557 190 559 193
rect 567 190 569 193
rect 577 190 579 193
rect 613 202 615 207
rect 623 202 625 207
rect 708 205 710 210
rect 718 205 720 210
rect 769 207 775 208
rect 769 203 770 207
rect 774 203 775 207
rect 769 202 775 203
rect 698 192 700 195
rect 708 192 710 195
rect 530 188 543 190
rect 549 188 559 190
rect 563 189 569 190
rect 489 184 495 185
rect 458 183 467 184
rect 390 176 391 180
rect 395 176 396 180
rect 390 175 396 176
rect 390 172 392 175
rect 371 165 373 169
rect 458 179 459 183
rect 463 179 467 183
rect 483 180 485 184
rect 458 178 467 179
rect 465 175 467 178
rect 475 175 477 180
rect 483 178 487 180
rect 485 175 487 178
rect 492 175 494 184
rect 533 180 535 188
rect 549 184 551 188
rect 563 185 564 189
rect 568 185 569 189
rect 563 184 569 185
rect 573 189 579 190
rect 573 185 574 189
rect 578 185 579 189
rect 573 184 579 185
rect 603 189 605 192
rect 613 189 615 192
rect 603 188 609 189
rect 603 184 604 188
rect 608 184 609 188
rect 613 186 617 189
rect 542 183 551 184
rect 449 168 451 171
rect 449 166 454 168
rect 240 156 242 161
rect 247 156 249 161
rect 207 154 232 156
rect 286 156 288 161
rect 293 156 295 161
rect 383 158 385 163
rect 390 158 392 163
rect 452 158 454 166
rect 465 162 467 166
rect 475 158 477 166
rect 542 179 543 183
rect 547 179 551 183
rect 567 180 569 184
rect 542 178 551 179
rect 549 175 551 178
rect 559 175 561 180
rect 567 178 571 180
rect 569 175 571 178
rect 576 175 578 184
rect 603 183 609 184
rect 603 175 605 183
rect 533 168 535 171
rect 533 166 538 168
rect 485 158 487 163
rect 492 158 494 163
rect 452 156 477 158
rect 536 158 538 166
rect 549 162 551 166
rect 559 158 561 166
rect 615 172 617 186
rect 623 181 625 192
rect 698 191 704 192
rect 698 187 699 191
rect 703 187 704 191
rect 708 189 712 192
rect 698 186 704 187
rect 622 180 628 181
rect 622 176 623 180
rect 627 176 628 180
rect 698 178 700 186
rect 622 175 628 176
rect 622 172 624 175
rect 710 175 712 189
rect 718 184 720 195
rect 773 193 775 202
rect 820 223 822 227
rect 868 223 870 227
rect 800 214 802 218
rect 810 214 812 218
rect 853 207 859 208
rect 853 203 854 207
rect 858 203 859 207
rect 853 202 859 203
rect 784 193 786 196
rect 800 193 802 196
rect 810 193 812 196
rect 820 193 822 196
rect 773 191 786 193
rect 792 191 802 193
rect 806 192 812 193
rect 717 183 723 184
rect 776 183 778 191
rect 792 187 794 191
rect 806 188 807 192
rect 811 188 812 192
rect 806 187 812 188
rect 816 192 822 193
rect 816 188 817 192
rect 821 188 822 192
rect 857 193 859 202
rect 904 223 906 227
rect 884 214 886 218
rect 894 214 896 218
rect 940 215 946 216
rect 930 207 932 212
rect 940 211 941 215
rect 945 211 946 215
rect 940 210 946 211
rect 868 193 870 196
rect 884 193 886 196
rect 894 193 896 196
rect 904 193 906 196
rect 940 205 942 210
rect 950 205 952 210
rect 1118 206 1120 224
rect 1157 206 1159 221
rect 1178 206 1180 221
rect 1211 206 1213 221
rect 1232 206 1234 221
rect 1267 206 1269 221
rect 1288 206 1290 221
rect 1321 206 1323 221
rect 1342 206 1344 221
rect 1158 202 1159 206
rect 1179 202 1180 206
rect 1212 202 1213 206
rect 1233 202 1234 206
rect 1268 202 1269 206
rect 1289 202 1290 206
rect 1322 202 1323 206
rect 1343 202 1344 206
rect 857 191 870 193
rect 876 191 886 193
rect 890 192 896 193
rect 816 187 822 188
rect 785 186 794 187
rect 717 179 718 183
rect 722 179 723 183
rect 717 178 723 179
rect 717 175 719 178
rect 603 165 605 169
rect 698 168 700 172
rect 785 182 786 186
rect 790 182 794 186
rect 810 183 812 187
rect 785 181 794 182
rect 792 178 794 181
rect 802 178 804 183
rect 810 181 814 183
rect 812 178 814 181
rect 819 178 821 187
rect 860 183 862 191
rect 876 187 878 191
rect 890 188 891 192
rect 895 188 896 192
rect 890 187 896 188
rect 900 192 906 193
rect 900 188 901 192
rect 905 188 906 192
rect 900 187 906 188
rect 930 192 932 195
rect 940 192 942 195
rect 930 191 936 192
rect 930 187 931 191
rect 935 187 936 191
rect 940 189 944 192
rect 869 186 878 187
rect 776 171 778 174
rect 776 169 781 171
rect 569 158 571 163
rect 576 158 578 163
rect 536 156 561 158
rect 615 158 617 163
rect 622 158 624 163
rect 710 161 712 166
rect 717 161 719 166
rect 779 161 781 169
rect 792 165 794 169
rect 802 161 804 169
rect 869 182 870 186
rect 874 182 878 186
rect 894 183 896 187
rect 869 181 878 182
rect 876 178 878 181
rect 886 178 888 183
rect 894 181 898 183
rect 896 178 898 181
rect 903 178 905 187
rect 930 186 936 187
rect 930 178 932 186
rect 860 171 862 174
rect 860 169 865 171
rect 812 161 814 166
rect 819 161 821 166
rect 779 159 804 161
rect 863 161 865 169
rect 876 165 878 169
rect 886 161 888 169
rect 942 175 944 189
rect 950 184 952 195
rect 1118 190 1120 202
rect 1157 190 1159 202
rect 1178 190 1180 202
rect 1211 190 1213 202
rect 1232 190 1234 202
rect 1267 190 1269 202
rect 1288 190 1290 202
rect 1321 190 1323 202
rect 1342 190 1344 202
rect 949 183 955 184
rect 949 179 950 183
rect 954 179 955 183
rect 949 178 955 179
rect 1118 178 1120 184
rect 1157 178 1159 184
rect 1178 178 1180 184
rect 1211 178 1213 184
rect 1232 178 1234 184
rect 1267 178 1269 184
rect 1288 178 1290 184
rect 1321 178 1323 184
rect 1342 178 1344 184
rect 949 175 951 178
rect 930 168 932 172
rect 896 161 898 166
rect 903 161 905 166
rect 863 159 888 161
rect 942 161 944 166
rect 949 161 951 166
rect 135 139 137 143
rect 145 139 147 143
rect 155 139 157 143
rect 464 141 466 145
rect 474 141 476 145
rect 484 141 486 145
rect 791 144 793 148
rect 801 144 803 148
rect 811 144 813 148
rect 1041 147 1043 149
rect 1113 147 1115 153
rect 1152 147 1154 153
rect 1173 147 1175 153
rect 1206 147 1208 153
rect 1227 147 1229 153
rect 1262 147 1264 153
rect 1283 147 1285 153
rect 1316 147 1318 153
rect 1337 147 1339 153
rect 135 125 137 133
rect 131 124 137 125
rect 145 124 147 133
rect 155 124 157 133
rect 464 127 466 135
rect 131 120 132 124
rect 136 120 137 124
rect 151 123 157 124
rect 131 119 137 120
rect 135 106 137 119
rect 145 117 147 120
rect 151 119 152 123
rect 156 119 157 123
rect 460 126 466 127
rect 474 126 476 135
rect 484 126 486 135
rect 791 130 793 138
rect 460 122 461 126
rect 465 122 466 126
rect 480 125 486 126
rect 460 121 466 122
rect 151 118 157 119
rect 141 116 147 117
rect 141 112 142 116
rect 146 112 147 116
rect 141 111 147 112
rect 142 106 144 111
rect 155 109 157 118
rect 464 108 466 121
rect 474 119 476 122
rect 480 121 481 125
rect 485 121 486 125
rect 787 129 793 130
rect 801 129 803 138
rect 811 129 813 138
rect 1041 130 1043 141
rect 787 125 788 129
rect 792 125 793 129
rect 807 128 813 129
rect 787 124 793 125
rect 480 120 486 121
rect 470 118 476 119
rect 470 114 471 118
rect 475 114 476 118
rect 470 113 476 114
rect 471 108 473 113
rect 484 111 486 120
rect 791 111 793 124
rect 801 122 803 125
rect 807 124 808 128
rect 812 124 813 128
rect 1113 129 1115 141
rect 1152 129 1154 141
rect 1173 129 1175 141
rect 1206 129 1208 141
rect 1227 129 1229 141
rect 1262 129 1264 141
rect 1283 129 1285 141
rect 1316 129 1318 141
rect 1337 129 1339 141
rect 807 123 813 124
rect 797 121 803 122
rect 797 117 798 121
rect 802 117 803 121
rect 797 116 803 117
rect 798 111 800 116
rect 811 114 813 123
rect 155 93 157 97
rect 484 95 486 99
rect 1041 108 1043 126
rect 1153 125 1154 129
rect 1174 125 1175 129
rect 1207 125 1208 129
rect 1228 125 1229 129
rect 1263 125 1264 129
rect 1284 125 1285 129
rect 1317 125 1318 129
rect 1338 125 1339 129
rect 1041 102 1043 105
rect 1113 107 1115 125
rect 1152 110 1154 125
rect 1173 110 1175 125
rect 1206 110 1208 125
rect 1227 110 1229 125
rect 1262 110 1264 125
rect 1283 110 1285 125
rect 1316 110 1318 125
rect 1337 110 1339 125
rect 811 98 813 102
rect 1113 101 1115 104
rect 1152 101 1154 104
rect 1173 101 1175 104
rect 1206 101 1208 104
rect 1227 101 1229 104
rect 1262 101 1264 104
rect 1283 101 1285 104
rect 1316 101 1318 104
rect 1337 101 1339 104
rect 135 84 137 88
rect 142 84 144 88
rect 464 86 466 90
rect 471 86 473 90
rect 791 89 793 93
rect 798 89 800 93
rect 1117 85 1119 88
rect 1156 85 1158 88
rect 1177 85 1179 88
rect 1210 85 1212 88
rect 1231 85 1233 88
rect 1266 85 1268 88
rect 1287 85 1289 88
rect 1320 85 1322 88
rect 1341 85 1343 88
rect 336 61 338 65
rect 346 63 348 68
rect 356 63 358 68
rect 429 61 431 65
rect 439 63 441 68
rect 449 63 451 68
rect 336 39 338 43
rect 346 39 348 50
rect 356 47 358 50
rect 356 46 362 47
rect 356 42 357 46
rect 361 42 362 46
rect 516 61 518 65
rect 526 63 528 68
rect 536 63 538 68
rect 1117 64 1119 82
rect 1156 64 1158 79
rect 1177 64 1179 79
rect 1210 64 1212 79
rect 1231 64 1233 79
rect 1266 64 1268 79
rect 1287 64 1289 79
rect 1320 64 1322 79
rect 1341 64 1343 79
rect 356 41 362 42
rect 336 38 342 39
rect 336 34 337 38
rect 341 34 342 38
rect 336 33 342 34
rect 346 38 352 39
rect 346 34 347 38
rect 351 34 352 38
rect 346 33 352 34
rect 336 28 338 33
rect 349 28 351 33
rect 356 28 358 41
rect 429 39 431 43
rect 439 39 441 50
rect 449 47 451 50
rect 449 46 455 47
rect 449 42 450 46
rect 454 42 455 46
rect 1157 60 1158 64
rect 1178 60 1179 64
rect 1211 60 1212 64
rect 1232 60 1233 64
rect 1267 60 1268 64
rect 1288 60 1289 64
rect 1321 60 1322 64
rect 1342 60 1343 64
rect 449 41 455 42
rect 429 38 435 39
rect 429 34 430 38
rect 434 34 435 38
rect 429 33 435 34
rect 439 38 445 39
rect 439 34 440 38
rect 444 34 445 38
rect 439 33 445 34
rect 429 28 431 33
rect 442 28 444 33
rect 449 28 451 41
rect 516 39 518 43
rect 526 39 528 50
rect 536 47 538 50
rect 1117 48 1119 60
rect 1156 48 1158 60
rect 1177 48 1179 60
rect 1210 48 1212 60
rect 1231 48 1233 60
rect 1266 48 1268 60
rect 1287 48 1289 60
rect 1320 48 1322 60
rect 1341 48 1343 60
rect 536 46 542 47
rect 536 42 537 46
rect 541 42 542 46
rect 536 41 542 42
rect 516 38 522 39
rect 516 34 517 38
rect 521 34 522 38
rect 516 33 522 34
rect 526 38 532 39
rect 526 34 527 38
rect 531 34 532 38
rect 526 33 532 34
rect 516 28 518 33
rect 529 28 531 33
rect 536 28 538 41
rect 1117 36 1119 42
rect 1156 36 1158 42
rect 1177 36 1179 42
rect 1210 36 1212 42
rect 1231 36 1233 42
rect 1266 36 1268 42
rect 1287 36 1289 42
rect 1320 36 1322 42
rect 1341 36 1343 42
rect 336 15 338 19
rect 349 12 351 17
rect 356 12 358 17
rect 429 15 431 19
rect 442 12 444 17
rect 449 12 451 17
rect 516 15 518 19
rect 529 12 531 17
rect 536 12 538 17
<< ndiffusion >>
rect 132 445 139 446
rect 132 441 134 445
rect 138 441 139 445
rect 132 436 139 441
rect 219 445 226 446
rect 219 441 221 445
rect 225 441 226 445
rect 114 435 121 436
rect 114 431 115 435
rect 119 431 121 435
rect 114 430 121 431
rect 116 425 121 430
rect 123 425 128 436
rect 130 434 139 436
rect 219 436 226 441
rect 312 445 319 446
rect 312 441 314 445
rect 318 441 319 445
rect 201 435 208 436
rect 130 425 141 434
rect 143 433 150 434
rect 143 429 145 433
rect 149 429 150 433
rect 201 431 202 435
rect 206 431 208 435
rect 201 430 208 431
rect 143 428 150 429
rect 143 425 148 428
rect 203 425 208 430
rect 210 425 215 436
rect 217 434 226 436
rect 312 436 319 441
rect 545 447 552 448
rect 545 443 546 447
rect 550 443 552 447
rect 294 435 301 436
rect 217 425 228 434
rect 230 433 237 434
rect 230 429 232 433
rect 236 429 237 433
rect 294 431 295 435
rect 299 431 301 435
rect 294 430 301 431
rect 230 428 237 429
rect 230 425 235 428
rect 296 425 301 430
rect 303 425 308 436
rect 310 434 319 436
rect 545 438 552 443
rect 638 447 645 448
rect 638 443 639 447
rect 643 443 645 447
rect 545 436 554 438
rect 534 435 541 436
rect 310 425 321 434
rect 323 433 330 434
rect 323 429 325 433
rect 329 429 330 433
rect 534 431 535 435
rect 539 431 541 435
rect 534 430 541 431
rect 323 428 330 429
rect 323 425 328 428
rect 536 427 541 430
rect 543 427 554 436
rect 556 427 561 438
rect 563 437 570 438
rect 563 433 565 437
rect 569 433 570 437
rect 638 438 645 443
rect 725 447 732 448
rect 725 443 726 447
rect 730 443 732 447
rect 638 436 647 438
rect 563 432 570 433
rect 627 435 634 436
rect 563 427 568 432
rect 627 431 628 435
rect 632 431 634 435
rect 627 430 634 431
rect 629 427 634 430
rect 636 427 647 436
rect 649 427 654 438
rect 656 437 663 438
rect 656 433 658 437
rect 662 433 663 437
rect 725 438 732 443
rect 725 436 734 438
rect 656 432 663 433
rect 714 435 721 436
rect 656 427 661 432
rect 714 431 715 435
rect 719 431 721 435
rect 714 430 721 431
rect 716 427 721 430
rect 723 427 734 436
rect 736 427 741 438
rect 743 437 750 438
rect 743 433 745 437
rect 749 433 750 437
rect 743 432 750 433
rect 743 427 748 432
rect 1031 392 1042 395
rect 1044 392 1061 395
rect 1143 396 1153 397
rect 1103 391 1114 394
rect 1116 391 1133 394
rect 1143 392 1145 396
rect 1149 392 1153 396
rect 1143 391 1153 392
rect 1155 391 1174 397
rect 1176 396 1184 397
rect 1176 392 1179 396
rect 1183 392 1184 396
rect 1176 391 1184 392
rect 1197 396 1207 397
rect 1197 392 1199 396
rect 1203 392 1207 396
rect 1197 391 1207 392
rect 1209 391 1228 397
rect 1230 396 1238 397
rect 1230 392 1233 396
rect 1237 392 1238 396
rect 1230 391 1238 392
rect 1253 396 1263 397
rect 1253 392 1255 396
rect 1259 392 1263 396
rect 1253 391 1263 392
rect 1265 391 1284 397
rect 1286 396 1294 397
rect 1286 392 1289 396
rect 1293 392 1294 396
rect 1286 391 1294 392
rect 1307 396 1317 397
rect 1307 392 1309 396
rect 1313 392 1317 396
rect 1307 391 1317 392
rect 1319 391 1338 397
rect 1340 396 1348 397
rect 1340 392 1343 396
rect 1347 392 1348 396
rect 1340 391 1348 392
rect 36 318 43 319
rect 36 314 37 318
rect 41 314 43 318
rect 36 313 43 314
rect 45 316 53 319
rect 114 323 121 324
rect 114 319 115 323
rect 119 319 121 323
rect 114 318 121 319
rect 45 313 55 316
rect 47 307 55 313
rect 57 307 62 316
rect 64 315 71 316
rect 116 315 121 318
rect 123 319 128 324
rect 198 323 205 324
rect 198 319 199 323
rect 203 319 205 323
rect 123 315 137 319
rect 64 311 66 315
rect 70 311 71 315
rect 64 310 71 311
rect 128 311 129 315
rect 133 311 137 315
rect 128 310 137 311
rect 139 318 147 319
rect 139 314 141 318
rect 145 314 147 318
rect 139 310 147 314
rect 149 316 157 319
rect 149 312 151 316
rect 155 312 157 316
rect 149 310 157 312
rect 64 307 69 310
rect 47 306 53 307
rect 47 302 48 306
rect 52 302 53 306
rect 47 301 53 302
rect 152 307 157 310
rect 159 307 164 319
rect 166 307 174 319
rect 198 318 205 319
rect 200 315 205 318
rect 207 319 212 324
rect 207 315 221 319
rect 212 311 213 315
rect 217 311 221 315
rect 212 310 221 311
rect 223 318 231 319
rect 223 314 225 318
rect 229 314 231 318
rect 223 310 231 314
rect 233 316 241 319
rect 233 312 235 316
rect 239 312 241 316
rect 233 310 241 312
rect 168 306 174 307
rect 168 302 169 306
rect 173 302 174 306
rect 168 301 174 302
rect 236 307 241 310
rect 243 307 248 319
rect 250 307 258 319
rect 268 318 275 319
rect 268 314 269 318
rect 273 314 275 318
rect 268 313 275 314
rect 277 316 285 319
rect 365 320 372 321
rect 365 316 366 320
rect 370 316 372 320
rect 277 313 287 316
rect 279 307 287 313
rect 289 307 294 316
rect 296 315 303 316
rect 365 315 372 316
rect 374 318 382 321
rect 443 325 450 326
rect 443 321 444 325
rect 448 321 450 325
rect 443 320 450 321
rect 374 315 384 318
rect 296 311 298 315
rect 302 311 303 315
rect 296 310 303 311
rect 296 307 301 310
rect 376 309 384 315
rect 386 309 391 318
rect 393 317 400 318
rect 445 317 450 320
rect 452 321 457 326
rect 527 325 534 326
rect 527 321 528 325
rect 532 321 534 325
rect 452 317 466 321
rect 393 313 395 317
rect 399 313 400 317
rect 393 312 400 313
rect 457 313 458 317
rect 462 313 466 317
rect 457 312 466 313
rect 468 320 476 321
rect 468 316 470 320
rect 474 316 476 320
rect 468 312 476 316
rect 478 318 486 321
rect 478 314 480 318
rect 484 314 486 318
rect 478 312 486 314
rect 393 309 398 312
rect 252 306 258 307
rect 252 302 253 306
rect 257 302 258 306
rect 252 301 258 302
rect 279 306 285 307
rect 279 302 280 306
rect 284 302 285 306
rect 376 308 382 309
rect 376 304 377 308
rect 381 304 382 308
rect 376 303 382 304
rect 481 309 486 312
rect 488 309 493 321
rect 495 309 503 321
rect 527 320 534 321
rect 529 317 534 320
rect 536 321 541 326
rect 536 317 550 321
rect 541 313 542 317
rect 546 313 550 317
rect 541 312 550 313
rect 552 320 560 321
rect 552 316 554 320
rect 558 316 560 320
rect 552 312 560 316
rect 562 318 570 321
rect 562 314 564 318
rect 568 314 570 318
rect 562 312 570 314
rect 497 308 503 309
rect 497 304 498 308
rect 502 304 503 308
rect 497 303 503 304
rect 565 309 570 312
rect 572 309 577 321
rect 579 309 587 321
rect 597 320 604 321
rect 597 316 598 320
rect 602 316 604 320
rect 597 315 604 316
rect 606 318 614 321
rect 692 323 699 324
rect 692 319 693 323
rect 697 319 699 323
rect 692 318 699 319
rect 701 321 709 324
rect 1107 369 1118 372
rect 1120 369 1137 372
rect 1147 371 1157 372
rect 1147 367 1149 371
rect 1153 367 1157 371
rect 1147 366 1157 367
rect 1159 366 1178 372
rect 1180 371 1188 372
rect 1180 367 1183 371
rect 1187 367 1188 371
rect 1180 366 1188 367
rect 1201 371 1211 372
rect 1201 367 1203 371
rect 1207 367 1211 371
rect 1201 366 1211 367
rect 1213 366 1232 372
rect 1234 371 1242 372
rect 1234 367 1237 371
rect 1241 367 1242 371
rect 1234 366 1242 367
rect 1257 371 1267 372
rect 1257 367 1259 371
rect 1263 367 1267 371
rect 1257 366 1267 367
rect 1269 366 1288 372
rect 1290 371 1298 372
rect 1290 367 1293 371
rect 1297 367 1298 371
rect 1290 366 1298 367
rect 1311 371 1321 372
rect 1311 367 1313 371
rect 1317 367 1321 371
rect 1311 366 1321 367
rect 1323 366 1342 372
rect 1344 371 1352 372
rect 1344 367 1347 371
rect 1351 367 1352 371
rect 1344 366 1352 367
rect 770 328 777 329
rect 770 324 771 328
rect 775 324 777 328
rect 770 323 777 324
rect 701 318 711 321
rect 606 315 616 318
rect 608 309 616 315
rect 618 309 623 318
rect 625 317 632 318
rect 625 313 627 317
rect 631 313 632 317
rect 625 312 632 313
rect 703 312 711 318
rect 713 312 718 321
rect 720 320 727 321
rect 772 320 777 323
rect 779 324 784 329
rect 854 328 861 329
rect 854 324 855 328
rect 859 324 861 328
rect 779 320 793 324
rect 720 316 722 320
rect 726 316 727 320
rect 720 315 727 316
rect 784 316 785 320
rect 789 316 793 320
rect 784 315 793 316
rect 795 323 803 324
rect 795 319 797 323
rect 801 319 803 323
rect 795 315 803 319
rect 805 321 813 324
rect 805 317 807 321
rect 811 317 813 321
rect 805 315 813 317
rect 720 312 725 315
rect 625 309 630 312
rect 581 308 587 309
rect 581 304 582 308
rect 586 304 587 308
rect 581 303 587 304
rect 608 308 614 309
rect 608 304 609 308
rect 613 304 614 308
rect 703 311 709 312
rect 703 307 704 311
rect 708 307 709 311
rect 703 306 709 307
rect 808 312 813 315
rect 815 312 820 324
rect 822 312 830 324
rect 854 323 861 324
rect 856 320 861 323
rect 863 324 868 329
rect 863 320 877 324
rect 868 316 869 320
rect 873 316 877 320
rect 868 315 877 316
rect 879 323 887 324
rect 879 319 881 323
rect 885 319 887 323
rect 879 315 887 319
rect 889 321 897 324
rect 889 317 891 321
rect 895 317 897 321
rect 889 315 897 317
rect 824 311 830 312
rect 824 307 825 311
rect 829 307 830 311
rect 824 306 830 307
rect 892 312 897 315
rect 899 312 904 324
rect 906 312 914 324
rect 924 323 931 324
rect 924 319 925 323
rect 929 319 931 323
rect 924 318 931 319
rect 933 321 941 324
rect 933 318 943 321
rect 935 312 943 318
rect 945 312 950 321
rect 952 320 959 321
rect 952 316 954 320
rect 958 316 959 320
rect 952 315 959 316
rect 952 312 957 315
rect 908 311 914 312
rect 908 307 909 311
rect 913 307 914 311
rect 908 306 914 307
rect 935 311 941 312
rect 935 307 936 311
rect 940 307 941 311
rect 935 306 941 307
rect 608 303 614 304
rect 279 301 285 302
rect 785 289 792 290
rect 458 286 465 287
rect 129 284 136 285
rect 129 280 130 284
rect 134 280 136 284
rect 129 279 136 280
rect 138 284 146 285
rect 138 280 140 284
rect 144 280 146 284
rect 138 279 146 280
rect 148 284 156 285
rect 148 280 150 284
rect 154 280 156 284
rect 148 279 156 280
rect 158 284 165 285
rect 158 280 160 284
rect 164 280 165 284
rect 458 282 459 286
rect 463 282 465 286
rect 458 281 465 282
rect 467 286 475 287
rect 467 282 469 286
rect 473 282 475 286
rect 467 281 475 282
rect 477 286 485 287
rect 477 282 479 286
rect 483 282 485 286
rect 477 281 485 282
rect 487 286 494 287
rect 487 282 489 286
rect 493 282 494 286
rect 785 285 786 289
rect 790 285 792 289
rect 785 284 792 285
rect 794 289 802 290
rect 794 285 796 289
rect 800 285 802 289
rect 794 284 802 285
rect 804 289 812 290
rect 804 285 806 289
rect 810 285 812 289
rect 804 284 812 285
rect 814 289 821 290
rect 814 285 816 289
rect 820 285 821 289
rect 814 284 821 285
rect 487 281 494 282
rect 158 279 165 280
rect 1031 247 1042 250
rect 1044 247 1061 250
rect 1143 251 1153 252
rect 1103 246 1114 249
rect 1116 246 1133 249
rect 1143 247 1145 251
rect 1149 247 1153 251
rect 1143 246 1153 247
rect 1155 246 1174 252
rect 1176 251 1184 252
rect 1176 247 1179 251
rect 1183 247 1184 251
rect 1176 246 1184 247
rect 1197 251 1207 252
rect 1197 247 1199 251
rect 1203 247 1207 251
rect 1197 246 1207 247
rect 1209 246 1228 252
rect 1230 251 1238 252
rect 1230 247 1233 251
rect 1237 247 1238 251
rect 1230 246 1238 247
rect 1253 251 1263 252
rect 1253 247 1255 251
rect 1259 247 1263 251
rect 1253 246 1263 247
rect 1265 246 1284 252
rect 1286 251 1294 252
rect 1286 247 1289 251
rect 1293 247 1294 251
rect 1286 246 1294 247
rect 1307 251 1317 252
rect 1307 247 1309 251
rect 1313 247 1317 251
rect 1307 246 1317 247
rect 1319 246 1338 252
rect 1340 251 1348 252
rect 1340 247 1343 251
rect 1347 247 1348 251
rect 1340 246 1348 247
rect 35 172 42 173
rect 35 168 36 172
rect 40 168 42 172
rect 35 167 42 168
rect 44 170 52 173
rect 113 177 120 178
rect 113 173 114 177
rect 118 173 120 177
rect 113 172 120 173
rect 44 167 54 170
rect 46 161 54 167
rect 56 161 61 170
rect 63 169 70 170
rect 115 169 120 172
rect 122 173 127 178
rect 197 177 204 178
rect 197 173 198 177
rect 202 173 204 177
rect 122 169 136 173
rect 63 165 65 169
rect 69 165 70 169
rect 63 164 70 165
rect 127 165 128 169
rect 132 165 136 169
rect 127 164 136 165
rect 138 172 146 173
rect 138 168 140 172
rect 144 168 146 172
rect 138 164 146 168
rect 148 170 156 173
rect 148 166 150 170
rect 154 166 156 170
rect 148 164 156 166
rect 63 161 68 164
rect 46 160 52 161
rect 46 156 47 160
rect 51 156 52 160
rect 46 155 52 156
rect 151 161 156 164
rect 158 161 163 173
rect 165 161 173 173
rect 197 172 204 173
rect 199 169 204 172
rect 206 173 211 178
rect 206 169 220 173
rect 211 165 212 169
rect 216 165 220 169
rect 211 164 220 165
rect 222 172 230 173
rect 222 168 224 172
rect 228 168 230 172
rect 222 164 230 168
rect 232 170 240 173
rect 232 166 234 170
rect 238 166 240 170
rect 232 164 240 166
rect 167 160 173 161
rect 167 156 168 160
rect 172 156 173 160
rect 167 155 173 156
rect 235 161 240 164
rect 242 161 247 173
rect 249 161 257 173
rect 267 172 274 173
rect 267 168 268 172
rect 272 168 274 172
rect 267 167 274 168
rect 276 170 284 173
rect 364 174 371 175
rect 364 170 365 174
rect 369 170 371 174
rect 276 167 286 170
rect 278 161 286 167
rect 288 161 293 170
rect 295 169 302 170
rect 364 169 371 170
rect 373 172 381 175
rect 442 179 449 180
rect 442 175 443 179
rect 447 175 449 179
rect 442 174 449 175
rect 373 169 383 172
rect 295 165 297 169
rect 301 165 302 169
rect 295 164 302 165
rect 295 161 300 164
rect 375 163 383 169
rect 385 163 390 172
rect 392 171 399 172
rect 444 171 449 174
rect 451 175 456 180
rect 526 179 533 180
rect 526 175 527 179
rect 531 175 533 179
rect 451 171 465 175
rect 392 167 394 171
rect 398 167 399 171
rect 392 166 399 167
rect 456 167 457 171
rect 461 167 465 171
rect 456 166 465 167
rect 467 174 475 175
rect 467 170 469 174
rect 473 170 475 174
rect 467 166 475 170
rect 477 172 485 175
rect 477 168 479 172
rect 483 168 485 172
rect 477 166 485 168
rect 392 163 397 166
rect 251 160 257 161
rect 251 156 252 160
rect 256 156 257 160
rect 251 155 257 156
rect 278 160 284 161
rect 278 156 279 160
rect 283 156 284 160
rect 375 162 381 163
rect 375 158 376 162
rect 380 158 381 162
rect 375 157 381 158
rect 480 163 485 166
rect 487 163 492 175
rect 494 163 502 175
rect 526 174 533 175
rect 528 171 533 174
rect 535 175 540 180
rect 535 171 549 175
rect 540 167 541 171
rect 545 167 549 171
rect 540 166 549 167
rect 551 174 559 175
rect 551 170 553 174
rect 557 170 559 174
rect 551 166 559 170
rect 561 172 569 175
rect 561 168 563 172
rect 567 168 569 172
rect 561 166 569 168
rect 496 162 502 163
rect 496 158 497 162
rect 501 158 502 162
rect 496 157 502 158
rect 564 163 569 166
rect 571 163 576 175
rect 578 163 586 175
rect 596 174 603 175
rect 596 170 597 174
rect 601 170 603 174
rect 596 169 603 170
rect 605 172 613 175
rect 691 177 698 178
rect 691 173 692 177
rect 696 173 698 177
rect 691 172 698 173
rect 700 175 708 178
rect 1107 224 1118 227
rect 1120 224 1137 227
rect 1147 226 1157 227
rect 1147 222 1149 226
rect 1153 222 1157 226
rect 1147 221 1157 222
rect 1159 221 1178 227
rect 1180 226 1188 227
rect 1180 222 1183 226
rect 1187 222 1188 226
rect 1180 221 1188 222
rect 1201 226 1211 227
rect 1201 222 1203 226
rect 1207 222 1211 226
rect 1201 221 1211 222
rect 1213 221 1232 227
rect 1234 226 1242 227
rect 1234 222 1237 226
rect 1241 222 1242 226
rect 1234 221 1242 222
rect 1257 226 1267 227
rect 1257 222 1259 226
rect 1263 222 1267 226
rect 1257 221 1267 222
rect 1269 221 1288 227
rect 1290 226 1298 227
rect 1290 222 1293 226
rect 1297 222 1298 226
rect 1290 221 1298 222
rect 1311 226 1321 227
rect 1311 222 1313 226
rect 1317 222 1321 226
rect 1311 221 1321 222
rect 1323 221 1342 227
rect 1344 226 1352 227
rect 1344 222 1347 226
rect 1351 222 1352 226
rect 1344 221 1352 222
rect 769 182 776 183
rect 769 178 770 182
rect 774 178 776 182
rect 769 177 776 178
rect 700 172 710 175
rect 605 169 615 172
rect 607 163 615 169
rect 617 163 622 172
rect 624 171 631 172
rect 624 167 626 171
rect 630 167 631 171
rect 624 166 631 167
rect 702 166 710 172
rect 712 166 717 175
rect 719 174 726 175
rect 771 174 776 177
rect 778 178 783 183
rect 853 182 860 183
rect 853 178 854 182
rect 858 178 860 182
rect 778 174 792 178
rect 719 170 721 174
rect 725 170 726 174
rect 719 169 726 170
rect 783 170 784 174
rect 788 170 792 174
rect 783 169 792 170
rect 794 177 802 178
rect 794 173 796 177
rect 800 173 802 177
rect 794 169 802 173
rect 804 175 812 178
rect 804 171 806 175
rect 810 171 812 175
rect 804 169 812 171
rect 719 166 724 169
rect 624 163 629 166
rect 580 162 586 163
rect 580 158 581 162
rect 585 158 586 162
rect 580 157 586 158
rect 607 162 613 163
rect 607 158 608 162
rect 612 158 613 162
rect 702 165 708 166
rect 702 161 703 165
rect 707 161 708 165
rect 702 160 708 161
rect 807 166 812 169
rect 814 166 819 178
rect 821 166 829 178
rect 853 177 860 178
rect 855 174 860 177
rect 862 178 867 183
rect 862 174 876 178
rect 867 170 868 174
rect 872 170 876 174
rect 867 169 876 170
rect 878 177 886 178
rect 878 173 880 177
rect 884 173 886 177
rect 878 169 886 173
rect 888 175 896 178
rect 888 171 890 175
rect 894 171 896 175
rect 888 169 896 171
rect 823 165 829 166
rect 823 161 824 165
rect 828 161 829 165
rect 823 160 829 161
rect 891 166 896 169
rect 898 166 903 178
rect 905 166 913 178
rect 923 177 930 178
rect 923 173 924 177
rect 928 173 930 177
rect 923 172 930 173
rect 932 175 940 178
rect 932 172 942 175
rect 934 166 942 172
rect 944 166 949 175
rect 951 174 958 175
rect 951 170 953 174
rect 957 170 958 174
rect 951 169 958 170
rect 951 166 956 169
rect 907 165 913 166
rect 907 161 908 165
rect 912 161 913 165
rect 907 160 913 161
rect 934 165 940 166
rect 934 161 935 165
rect 939 161 940 165
rect 934 160 940 161
rect 607 157 613 158
rect 278 155 284 156
rect 784 143 791 144
rect 457 140 464 141
rect 128 138 135 139
rect 128 134 129 138
rect 133 134 135 138
rect 128 133 135 134
rect 137 138 145 139
rect 137 134 139 138
rect 143 134 145 138
rect 137 133 145 134
rect 147 138 155 139
rect 147 134 149 138
rect 153 134 155 138
rect 147 133 155 134
rect 157 138 164 139
rect 157 134 159 138
rect 163 134 164 138
rect 457 136 458 140
rect 462 136 464 140
rect 457 135 464 136
rect 466 140 474 141
rect 466 136 468 140
rect 472 136 474 140
rect 466 135 474 136
rect 476 140 484 141
rect 476 136 478 140
rect 482 136 484 140
rect 476 135 484 136
rect 486 140 493 141
rect 486 136 488 140
rect 492 136 493 140
rect 784 139 785 143
rect 789 139 791 143
rect 784 138 791 139
rect 793 143 801 144
rect 793 139 795 143
rect 799 139 801 143
rect 793 138 801 139
rect 803 143 811 144
rect 803 139 805 143
rect 809 139 811 143
rect 803 138 811 139
rect 813 143 820 144
rect 813 139 815 143
rect 819 139 820 143
rect 813 138 820 139
rect 486 135 493 136
rect 157 133 164 134
rect 1030 105 1041 108
rect 1043 105 1060 108
rect 1142 109 1152 110
rect 1102 104 1113 107
rect 1115 104 1132 107
rect 1142 105 1144 109
rect 1148 105 1152 109
rect 1142 104 1152 105
rect 1154 104 1173 110
rect 1175 109 1183 110
rect 1175 105 1178 109
rect 1182 105 1183 109
rect 1175 104 1183 105
rect 1196 109 1206 110
rect 1196 105 1198 109
rect 1202 105 1206 109
rect 1196 104 1206 105
rect 1208 104 1227 110
rect 1229 109 1237 110
rect 1229 105 1232 109
rect 1236 105 1237 109
rect 1229 104 1237 105
rect 1252 109 1262 110
rect 1252 105 1254 109
rect 1258 105 1262 109
rect 1252 104 1262 105
rect 1264 104 1283 110
rect 1285 109 1293 110
rect 1285 105 1288 109
rect 1292 105 1293 109
rect 1285 104 1293 105
rect 1306 109 1316 110
rect 1306 105 1308 109
rect 1312 105 1316 109
rect 1306 104 1316 105
rect 1318 104 1337 110
rect 1339 109 1347 110
rect 1339 105 1342 109
rect 1346 105 1347 109
rect 1339 104 1347 105
rect 1106 82 1117 85
rect 1119 82 1136 85
rect 1146 84 1156 85
rect 1146 80 1148 84
rect 1152 80 1156 84
rect 1146 79 1156 80
rect 1158 79 1177 85
rect 1179 84 1187 85
rect 1179 80 1182 84
rect 1186 80 1187 84
rect 1179 79 1187 80
rect 1200 84 1210 85
rect 1200 80 1202 84
rect 1206 80 1210 84
rect 1200 79 1210 80
rect 1212 79 1231 85
rect 1233 84 1241 85
rect 1233 80 1236 84
rect 1240 80 1241 84
rect 1233 79 1241 80
rect 1256 84 1266 85
rect 1256 80 1258 84
rect 1262 80 1266 84
rect 1256 79 1266 80
rect 1268 79 1287 85
rect 1289 84 1297 85
rect 1289 80 1292 84
rect 1296 80 1297 84
rect 1289 79 1297 80
rect 1310 84 1320 85
rect 1310 80 1312 84
rect 1316 80 1320 84
rect 1310 79 1320 80
rect 1322 79 1341 85
rect 1343 84 1351 85
rect 1343 80 1346 84
rect 1350 80 1351 84
rect 1343 79 1351 80
rect 331 25 336 28
rect 329 24 336 25
rect 329 20 330 24
rect 334 20 336 24
rect 329 19 336 20
rect 338 19 349 28
rect 340 17 349 19
rect 351 17 356 28
rect 358 23 363 28
rect 424 25 429 28
rect 422 24 429 25
rect 358 22 365 23
rect 358 18 360 22
rect 364 18 365 22
rect 422 20 423 24
rect 427 20 429 24
rect 422 19 429 20
rect 431 19 442 28
rect 358 17 365 18
rect 340 12 347 17
rect 433 17 442 19
rect 444 17 449 28
rect 451 23 456 28
rect 511 25 516 28
rect 509 24 516 25
rect 451 22 458 23
rect 451 18 453 22
rect 457 18 458 22
rect 509 20 510 24
rect 514 20 516 24
rect 509 19 516 20
rect 518 19 529 28
rect 451 17 458 18
rect 340 8 341 12
rect 345 8 347 12
rect 340 7 347 8
rect 433 12 440 17
rect 520 17 529 19
rect 531 17 536 28
rect 538 23 543 28
rect 538 22 545 23
rect 538 18 540 22
rect 544 18 545 22
rect 538 17 545 18
rect 433 8 434 12
rect 438 8 440 12
rect 433 7 440 8
rect 520 12 527 17
rect 520 8 521 12
rect 525 8 527 12
rect 520 7 527 8
<< pdiffusion >>
rect 1011 433 1042 434
rect 1011 429 1016 433
rect 1020 429 1042 433
rect 1011 428 1042 429
rect 1044 429 1060 434
rect 1066 429 1079 434
rect 1044 428 1079 429
rect 1099 433 1114 434
rect 1103 429 1114 433
rect 1099 428 1114 429
rect 1116 433 1136 434
rect 1116 429 1132 433
rect 1116 428 1136 429
rect 1143 433 1153 434
rect 1143 429 1145 433
rect 1149 429 1153 433
rect 1143 428 1153 429
rect 1155 433 1174 434
rect 1155 429 1162 433
rect 1166 429 1174 433
rect 1155 428 1174 429
rect 1176 433 1184 434
rect 1176 429 1179 433
rect 1183 429 1184 433
rect 1176 428 1184 429
rect 1197 433 1207 434
rect 1197 429 1199 433
rect 1203 429 1207 433
rect 1197 428 1207 429
rect 1209 433 1228 434
rect 1209 429 1216 433
rect 1220 429 1228 433
rect 1209 428 1228 429
rect 1230 433 1238 434
rect 1230 429 1233 433
rect 1237 429 1238 433
rect 1230 428 1238 429
rect 1253 433 1263 434
rect 1253 429 1255 433
rect 1259 429 1263 433
rect 1253 428 1263 429
rect 1265 433 1284 434
rect 1265 429 1272 433
rect 1276 429 1284 433
rect 1265 428 1284 429
rect 1286 433 1294 434
rect 1286 429 1289 433
rect 1293 429 1294 433
rect 1286 428 1294 429
rect 1307 433 1317 434
rect 1307 429 1309 433
rect 1313 429 1317 433
rect 1307 428 1317 429
rect 1319 433 1338 434
rect 1319 429 1326 433
rect 1330 429 1338 433
rect 1319 428 1338 429
rect 1340 433 1348 434
rect 1340 429 1343 433
rect 1347 429 1348 433
rect 1340 428 1348 429
rect 135 403 141 410
rect 114 395 121 403
rect 114 391 115 395
rect 119 391 121 395
rect 114 390 121 391
rect 123 402 131 403
rect 123 398 125 402
rect 129 398 131 402
rect 123 395 131 398
rect 123 391 125 395
rect 129 391 131 395
rect 123 390 131 391
rect 133 397 141 403
rect 133 393 135 397
rect 139 393 141 397
rect 133 392 141 393
rect 143 409 150 410
rect 143 405 145 409
rect 149 405 150 409
rect 143 402 150 405
rect 222 403 228 410
rect 143 398 145 402
rect 149 398 150 402
rect 143 397 150 398
rect 143 392 148 397
rect 201 395 208 403
rect 133 390 139 392
rect 201 391 202 395
rect 206 391 208 395
rect 201 390 208 391
rect 210 402 218 403
rect 210 398 212 402
rect 216 398 218 402
rect 210 395 218 398
rect 210 391 212 395
rect 216 391 218 395
rect 210 390 218 391
rect 220 397 228 403
rect 220 393 222 397
rect 226 393 228 397
rect 220 392 228 393
rect 230 409 237 410
rect 230 405 232 409
rect 236 405 237 409
rect 230 402 237 405
rect 534 411 541 412
rect 315 403 321 410
rect 230 398 232 402
rect 236 398 237 402
rect 230 397 237 398
rect 230 392 235 397
rect 294 395 301 403
rect 220 390 226 392
rect 294 391 295 395
rect 299 391 301 395
rect 294 390 301 391
rect 303 402 311 403
rect 303 398 305 402
rect 309 398 311 402
rect 303 395 311 398
rect 303 391 305 395
rect 309 391 311 395
rect 303 390 311 391
rect 313 397 321 403
rect 313 393 315 397
rect 319 393 321 397
rect 313 392 321 393
rect 323 409 330 410
rect 323 405 325 409
rect 329 405 330 409
rect 323 402 330 405
rect 323 398 325 402
rect 329 398 330 402
rect 534 407 535 411
rect 539 407 541 411
rect 534 404 541 407
rect 534 400 535 404
rect 539 400 541 404
rect 534 399 541 400
rect 323 397 330 398
rect 323 392 328 397
rect 536 394 541 399
rect 543 405 549 412
rect 627 411 634 412
rect 627 407 628 411
rect 632 407 634 411
rect 543 399 551 405
rect 543 395 545 399
rect 549 395 551 399
rect 543 394 551 395
rect 313 390 319 392
rect 545 392 551 394
rect 553 404 561 405
rect 553 400 555 404
rect 559 400 561 404
rect 553 397 561 400
rect 553 393 555 397
rect 559 393 561 397
rect 553 392 561 393
rect 563 397 570 405
rect 627 404 634 407
rect 627 400 628 404
rect 632 400 634 404
rect 627 399 634 400
rect 563 393 565 397
rect 569 393 570 397
rect 629 394 634 399
rect 636 405 642 412
rect 714 411 721 412
rect 714 407 715 411
rect 719 407 721 411
rect 636 399 644 405
rect 636 395 638 399
rect 642 395 644 399
rect 636 394 644 395
rect 563 392 570 393
rect 638 392 644 394
rect 646 404 654 405
rect 646 400 648 404
rect 652 400 654 404
rect 646 397 654 400
rect 646 393 648 397
rect 652 393 654 397
rect 646 392 654 393
rect 656 397 663 405
rect 714 404 721 407
rect 714 400 715 404
rect 719 400 721 404
rect 714 399 721 400
rect 656 393 658 397
rect 662 393 663 397
rect 716 394 721 399
rect 723 405 729 412
rect 723 399 731 405
rect 723 395 725 399
rect 729 395 731 399
rect 723 394 731 395
rect 656 392 663 393
rect 725 392 731 394
rect 733 404 741 405
rect 733 400 735 404
rect 739 400 741 404
rect 733 397 741 400
rect 733 393 735 397
rect 739 393 741 397
rect 733 392 741 393
rect 743 397 750 405
rect 743 393 745 397
rect 749 393 750 397
rect 743 392 750 393
rect 38 342 43 348
rect 36 341 43 342
rect 36 337 37 341
rect 41 337 43 341
rect 36 336 43 337
rect 45 346 51 348
rect 45 341 53 346
rect 45 337 47 341
rect 51 337 53 341
rect 45 336 53 337
rect 55 341 63 346
rect 55 337 57 341
rect 61 337 63 341
rect 55 336 63 337
rect 65 345 72 346
rect 65 341 67 345
rect 71 341 72 345
rect 124 343 129 364
rect 65 336 72 341
rect 122 342 129 343
rect 122 338 123 342
rect 127 338 129 342
rect 122 337 129 338
rect 131 363 143 364
rect 131 359 133 363
rect 137 359 143 363
rect 131 356 143 359
rect 131 352 133 356
rect 137 355 143 356
rect 160 355 165 364
rect 137 352 145 355
rect 131 337 145 352
rect 147 342 155 355
rect 147 338 149 342
rect 153 338 155 342
rect 147 337 155 338
rect 157 349 165 355
rect 157 345 159 349
rect 163 345 165 349
rect 157 337 165 345
rect 167 358 172 364
rect 167 357 174 358
rect 167 353 169 357
rect 173 353 174 357
rect 167 352 174 353
rect 167 337 172 352
rect 208 343 213 364
rect 206 342 213 343
rect 206 338 207 342
rect 211 338 213 342
rect 206 337 213 338
rect 215 363 227 364
rect 215 359 217 363
rect 221 359 227 363
rect 215 356 227 359
rect 215 352 217 356
rect 221 355 227 356
rect 244 355 249 364
rect 221 352 229 355
rect 215 337 229 352
rect 231 342 239 355
rect 231 338 233 342
rect 237 338 239 342
rect 231 337 239 338
rect 241 349 249 355
rect 241 345 243 349
rect 247 345 249 349
rect 241 337 249 345
rect 251 358 256 364
rect 251 357 258 358
rect 251 353 253 357
rect 257 353 258 357
rect 251 352 258 353
rect 251 337 256 352
rect 270 342 275 348
rect 268 341 275 342
rect 268 337 269 341
rect 273 337 275 341
rect 268 336 275 337
rect 277 346 283 348
rect 277 341 285 346
rect 277 337 279 341
rect 283 337 285 341
rect 277 336 285 337
rect 287 341 295 346
rect 287 337 289 341
rect 293 337 295 341
rect 287 336 295 337
rect 297 345 304 346
rect 297 341 299 345
rect 303 341 304 345
rect 367 344 372 350
rect 297 336 304 341
rect 365 343 372 344
rect 365 339 366 343
rect 370 339 372 343
rect 365 338 372 339
rect 374 348 380 350
rect 374 343 382 348
rect 374 339 376 343
rect 380 339 382 343
rect 374 338 382 339
rect 384 343 392 348
rect 384 339 386 343
rect 390 339 392 343
rect 384 338 392 339
rect 394 347 401 348
rect 394 343 396 347
rect 400 343 401 347
rect 453 345 458 366
rect 394 338 401 343
rect 451 344 458 345
rect 451 340 452 344
rect 456 340 458 344
rect 451 339 458 340
rect 460 365 472 366
rect 460 361 462 365
rect 466 361 472 365
rect 460 358 472 361
rect 460 354 462 358
rect 466 357 472 358
rect 489 357 494 366
rect 466 354 474 357
rect 460 339 474 354
rect 476 344 484 357
rect 476 340 478 344
rect 482 340 484 344
rect 476 339 484 340
rect 486 351 494 357
rect 486 347 488 351
rect 492 347 494 351
rect 486 339 494 347
rect 496 360 501 366
rect 496 359 503 360
rect 496 355 498 359
rect 502 355 503 359
rect 496 354 503 355
rect 496 339 501 354
rect 537 345 542 366
rect 535 344 542 345
rect 535 340 536 344
rect 540 340 542 344
rect 535 339 542 340
rect 544 365 556 366
rect 544 361 546 365
rect 550 361 556 365
rect 544 358 556 361
rect 544 354 546 358
rect 550 357 556 358
rect 573 357 578 366
rect 550 354 558 357
rect 544 339 558 354
rect 560 344 568 357
rect 560 340 562 344
rect 566 340 568 344
rect 560 339 568 340
rect 570 351 578 357
rect 570 347 572 351
rect 576 347 578 351
rect 570 339 578 347
rect 580 360 585 366
rect 580 359 587 360
rect 580 355 582 359
rect 586 355 587 359
rect 580 354 587 355
rect 580 339 585 354
rect 599 344 604 350
rect 597 343 604 344
rect 597 339 598 343
rect 602 339 604 343
rect 597 338 604 339
rect 606 348 612 350
rect 606 343 614 348
rect 606 339 608 343
rect 612 339 614 343
rect 606 338 614 339
rect 616 343 624 348
rect 616 339 618 343
rect 622 339 624 343
rect 616 338 624 339
rect 626 347 633 348
rect 694 347 699 353
rect 626 343 628 347
rect 632 343 633 347
rect 626 338 633 343
rect 692 346 699 347
rect 692 342 693 346
rect 697 342 699 346
rect 692 341 699 342
rect 701 351 707 353
rect 701 346 709 351
rect 701 342 703 346
rect 707 342 709 346
rect 701 341 709 342
rect 711 346 719 351
rect 711 342 713 346
rect 717 342 719 346
rect 711 341 719 342
rect 721 350 728 351
rect 721 346 723 350
rect 727 346 728 350
rect 780 348 785 369
rect 721 341 728 346
rect 778 347 785 348
rect 778 343 779 347
rect 783 343 785 347
rect 778 342 785 343
rect 787 368 799 369
rect 787 364 789 368
rect 793 364 799 368
rect 787 361 799 364
rect 787 357 789 361
rect 793 360 799 361
rect 816 360 821 369
rect 793 357 801 360
rect 787 342 801 357
rect 803 347 811 360
rect 803 343 805 347
rect 809 343 811 347
rect 803 342 811 343
rect 813 354 821 360
rect 813 350 815 354
rect 819 350 821 354
rect 813 342 821 350
rect 823 363 828 369
rect 823 362 830 363
rect 823 358 825 362
rect 829 358 830 362
rect 823 357 830 358
rect 823 342 828 357
rect 864 348 869 369
rect 862 347 869 348
rect 862 343 863 347
rect 867 343 869 347
rect 862 342 869 343
rect 871 368 883 369
rect 871 364 873 368
rect 877 364 883 368
rect 871 361 883 364
rect 871 357 873 361
rect 877 360 883 361
rect 900 360 905 369
rect 877 357 885 360
rect 871 342 885 357
rect 887 347 895 360
rect 887 343 889 347
rect 893 343 895 347
rect 887 342 895 343
rect 897 354 905 360
rect 897 350 899 354
rect 903 350 905 354
rect 897 342 905 350
rect 907 363 912 369
rect 907 362 914 363
rect 907 358 909 362
rect 913 358 914 362
rect 907 357 914 358
rect 907 342 912 357
rect 926 347 931 353
rect 924 346 931 347
rect 924 342 925 346
rect 929 342 931 346
rect 924 341 931 342
rect 933 351 939 353
rect 933 346 941 351
rect 933 342 935 346
rect 939 342 941 346
rect 933 341 941 342
rect 943 346 951 351
rect 943 342 945 346
rect 949 342 951 346
rect 943 341 951 342
rect 953 350 960 351
rect 953 346 955 350
rect 959 346 960 350
rect 953 341 960 346
rect 1103 334 1118 335
rect 1107 330 1118 334
rect 1103 329 1118 330
rect 1120 334 1140 335
rect 1120 330 1136 334
rect 1120 329 1140 330
rect 1147 334 1157 335
rect 1147 330 1149 334
rect 1153 330 1157 334
rect 1147 329 1157 330
rect 1159 334 1178 335
rect 1159 330 1166 334
rect 1170 330 1178 334
rect 1159 329 1178 330
rect 1180 334 1188 335
rect 1180 330 1183 334
rect 1187 330 1188 334
rect 1180 329 1188 330
rect 1201 334 1211 335
rect 1201 330 1203 334
rect 1207 330 1211 334
rect 1201 329 1211 330
rect 1213 334 1232 335
rect 1213 330 1220 334
rect 1224 330 1232 334
rect 1213 329 1232 330
rect 1234 334 1242 335
rect 1234 330 1237 334
rect 1241 330 1242 334
rect 1234 329 1242 330
rect 1257 334 1267 335
rect 1257 330 1259 334
rect 1263 330 1267 334
rect 1257 329 1267 330
rect 1269 334 1288 335
rect 1269 330 1276 334
rect 1280 330 1288 334
rect 1269 329 1288 330
rect 1290 334 1298 335
rect 1290 330 1293 334
rect 1297 330 1298 334
rect 1290 329 1298 330
rect 1311 334 1321 335
rect 1311 330 1313 334
rect 1317 330 1321 334
rect 1311 329 1321 330
rect 1323 334 1342 335
rect 1323 330 1330 334
rect 1334 330 1342 334
rect 1323 329 1342 330
rect 1344 334 1352 335
rect 1344 330 1347 334
rect 1351 330 1352 334
rect 1344 329 1352 330
rect 1011 288 1042 289
rect 1011 284 1016 288
rect 1020 284 1042 288
rect 148 252 156 255
rect 131 247 136 252
rect 129 246 136 247
rect 129 242 130 246
rect 134 242 136 246
rect 129 241 136 242
rect 131 234 136 241
rect 138 234 143 252
rect 145 243 156 252
rect 158 249 163 255
rect 1011 283 1042 284
rect 1044 284 1060 289
rect 1066 284 1079 289
rect 1044 283 1079 284
rect 1099 288 1114 289
rect 1103 284 1114 288
rect 1099 283 1114 284
rect 1116 288 1136 289
rect 1116 284 1132 288
rect 1116 283 1136 284
rect 1143 288 1153 289
rect 1143 284 1145 288
rect 1149 284 1153 288
rect 1143 283 1153 284
rect 1155 288 1174 289
rect 1155 284 1162 288
rect 1166 284 1174 288
rect 1155 283 1174 284
rect 1176 288 1184 289
rect 1176 284 1179 288
rect 1183 284 1184 288
rect 1176 283 1184 284
rect 1197 288 1207 289
rect 1197 284 1199 288
rect 1203 284 1207 288
rect 1197 283 1207 284
rect 1209 288 1228 289
rect 1209 284 1216 288
rect 1220 284 1228 288
rect 1209 283 1228 284
rect 1230 288 1238 289
rect 1230 284 1233 288
rect 1237 284 1238 288
rect 1230 283 1238 284
rect 1253 288 1263 289
rect 1253 284 1255 288
rect 1259 284 1263 288
rect 1253 283 1263 284
rect 1265 288 1284 289
rect 1265 284 1272 288
rect 1276 284 1284 288
rect 1265 283 1284 284
rect 1286 288 1294 289
rect 1286 284 1289 288
rect 1293 284 1294 288
rect 1286 283 1294 284
rect 1307 288 1317 289
rect 1307 284 1309 288
rect 1313 284 1317 288
rect 1307 283 1317 284
rect 1319 288 1338 289
rect 1319 284 1326 288
rect 1330 284 1338 288
rect 1319 283 1338 284
rect 1340 288 1348 289
rect 1340 284 1343 288
rect 1347 284 1348 288
rect 1340 283 1348 284
rect 804 257 812 260
rect 477 254 485 257
rect 460 249 465 254
rect 158 248 165 249
rect 158 244 160 248
rect 164 244 165 248
rect 158 243 165 244
rect 458 248 465 249
rect 458 244 459 248
rect 463 244 465 248
rect 458 243 465 244
rect 145 239 154 243
rect 145 235 148 239
rect 152 235 154 239
rect 145 234 154 235
rect 460 236 465 243
rect 467 236 472 254
rect 474 245 485 254
rect 487 251 492 257
rect 787 252 792 257
rect 785 251 792 252
rect 487 250 494 251
rect 487 246 489 250
rect 493 246 494 250
rect 785 247 786 251
rect 790 247 792 251
rect 785 246 792 247
rect 487 245 494 246
rect 474 241 483 245
rect 474 237 477 241
rect 481 237 483 241
rect 787 239 792 246
rect 794 239 799 257
rect 801 248 812 257
rect 814 254 819 260
rect 814 253 821 254
rect 814 249 816 253
rect 820 249 821 253
rect 814 248 821 249
rect 801 244 810 248
rect 801 240 804 244
rect 808 240 810 244
rect 801 239 810 240
rect 474 236 483 237
rect 37 196 42 202
rect 35 195 42 196
rect 35 191 36 195
rect 40 191 42 195
rect 35 190 42 191
rect 44 200 50 202
rect 44 195 52 200
rect 44 191 46 195
rect 50 191 52 195
rect 44 190 52 191
rect 54 195 62 200
rect 54 191 56 195
rect 60 191 62 195
rect 54 190 62 191
rect 64 199 71 200
rect 64 195 66 199
rect 70 195 71 199
rect 123 197 128 218
rect 64 190 71 195
rect 121 196 128 197
rect 121 192 122 196
rect 126 192 128 196
rect 121 191 128 192
rect 130 217 142 218
rect 130 213 132 217
rect 136 213 142 217
rect 130 210 142 213
rect 130 206 132 210
rect 136 209 142 210
rect 159 209 164 218
rect 136 206 144 209
rect 130 191 144 206
rect 146 196 154 209
rect 146 192 148 196
rect 152 192 154 196
rect 146 191 154 192
rect 156 203 164 209
rect 156 199 158 203
rect 162 199 164 203
rect 156 191 164 199
rect 166 212 171 218
rect 166 211 173 212
rect 166 207 168 211
rect 172 207 173 211
rect 166 206 173 207
rect 166 191 171 206
rect 207 197 212 218
rect 205 196 212 197
rect 205 192 206 196
rect 210 192 212 196
rect 205 191 212 192
rect 214 217 226 218
rect 214 213 216 217
rect 220 213 226 217
rect 214 210 226 213
rect 214 206 216 210
rect 220 209 226 210
rect 243 209 248 218
rect 220 206 228 209
rect 214 191 228 206
rect 230 196 238 209
rect 230 192 232 196
rect 236 192 238 196
rect 230 191 238 192
rect 240 203 248 209
rect 240 199 242 203
rect 246 199 248 203
rect 240 191 248 199
rect 250 212 255 218
rect 250 211 257 212
rect 250 207 252 211
rect 256 207 257 211
rect 250 206 257 207
rect 250 191 255 206
rect 269 196 274 202
rect 267 195 274 196
rect 267 191 268 195
rect 272 191 274 195
rect 267 190 274 191
rect 276 200 282 202
rect 276 195 284 200
rect 276 191 278 195
rect 282 191 284 195
rect 276 190 284 191
rect 286 195 294 200
rect 286 191 288 195
rect 292 191 294 195
rect 286 190 294 191
rect 296 199 303 200
rect 296 195 298 199
rect 302 195 303 199
rect 366 198 371 204
rect 296 190 303 195
rect 364 197 371 198
rect 364 193 365 197
rect 369 193 371 197
rect 364 192 371 193
rect 373 202 379 204
rect 373 197 381 202
rect 373 193 375 197
rect 379 193 381 197
rect 373 192 381 193
rect 383 197 391 202
rect 383 193 385 197
rect 389 193 391 197
rect 383 192 391 193
rect 393 201 400 202
rect 393 197 395 201
rect 399 197 400 201
rect 452 199 457 220
rect 393 192 400 197
rect 450 198 457 199
rect 450 194 451 198
rect 455 194 457 198
rect 450 193 457 194
rect 459 219 471 220
rect 459 215 461 219
rect 465 215 471 219
rect 459 212 471 215
rect 459 208 461 212
rect 465 211 471 212
rect 488 211 493 220
rect 465 208 473 211
rect 459 193 473 208
rect 475 198 483 211
rect 475 194 477 198
rect 481 194 483 198
rect 475 193 483 194
rect 485 205 493 211
rect 485 201 487 205
rect 491 201 493 205
rect 485 193 493 201
rect 495 214 500 220
rect 495 213 502 214
rect 495 209 497 213
rect 501 209 502 213
rect 495 208 502 209
rect 495 193 500 208
rect 536 199 541 220
rect 534 198 541 199
rect 534 194 535 198
rect 539 194 541 198
rect 534 193 541 194
rect 543 219 555 220
rect 543 215 545 219
rect 549 215 555 219
rect 543 212 555 215
rect 543 208 545 212
rect 549 211 555 212
rect 572 211 577 220
rect 549 208 557 211
rect 543 193 557 208
rect 559 198 567 211
rect 559 194 561 198
rect 565 194 567 198
rect 559 193 567 194
rect 569 205 577 211
rect 569 201 571 205
rect 575 201 577 205
rect 569 193 577 201
rect 579 214 584 220
rect 579 213 586 214
rect 579 209 581 213
rect 585 209 586 213
rect 579 208 586 209
rect 579 193 584 208
rect 598 198 603 204
rect 596 197 603 198
rect 596 193 597 197
rect 601 193 603 197
rect 596 192 603 193
rect 605 202 611 204
rect 605 197 613 202
rect 605 193 607 197
rect 611 193 613 197
rect 605 192 613 193
rect 615 197 623 202
rect 615 193 617 197
rect 621 193 623 197
rect 615 192 623 193
rect 625 201 632 202
rect 693 201 698 207
rect 625 197 627 201
rect 631 197 632 201
rect 625 192 632 197
rect 691 200 698 201
rect 691 196 692 200
rect 696 196 698 200
rect 691 195 698 196
rect 700 205 706 207
rect 700 200 708 205
rect 700 196 702 200
rect 706 196 708 200
rect 700 195 708 196
rect 710 200 718 205
rect 710 196 712 200
rect 716 196 718 200
rect 710 195 718 196
rect 720 204 727 205
rect 720 200 722 204
rect 726 200 727 204
rect 779 202 784 223
rect 720 195 727 200
rect 777 201 784 202
rect 777 197 778 201
rect 782 197 784 201
rect 777 196 784 197
rect 786 222 798 223
rect 786 218 788 222
rect 792 218 798 222
rect 786 215 798 218
rect 786 211 788 215
rect 792 214 798 215
rect 815 214 820 223
rect 792 211 800 214
rect 786 196 800 211
rect 802 201 810 214
rect 802 197 804 201
rect 808 197 810 201
rect 802 196 810 197
rect 812 208 820 214
rect 812 204 814 208
rect 818 204 820 208
rect 812 196 820 204
rect 822 217 827 223
rect 822 216 829 217
rect 822 212 824 216
rect 828 212 829 216
rect 822 211 829 212
rect 822 196 827 211
rect 863 202 868 223
rect 861 201 868 202
rect 861 197 862 201
rect 866 197 868 201
rect 861 196 868 197
rect 870 222 882 223
rect 870 218 872 222
rect 876 218 882 222
rect 870 215 882 218
rect 870 211 872 215
rect 876 214 882 215
rect 899 214 904 223
rect 876 211 884 214
rect 870 196 884 211
rect 886 201 894 214
rect 886 197 888 201
rect 892 197 894 201
rect 886 196 894 197
rect 896 208 904 214
rect 896 204 898 208
rect 902 204 904 208
rect 896 196 904 204
rect 906 217 911 223
rect 906 216 913 217
rect 906 212 908 216
rect 912 212 913 216
rect 906 211 913 212
rect 906 196 911 211
rect 925 201 930 207
rect 923 200 930 201
rect 923 196 924 200
rect 928 196 930 200
rect 923 195 930 196
rect 932 205 938 207
rect 932 200 940 205
rect 932 196 934 200
rect 938 196 940 200
rect 932 195 940 196
rect 942 200 950 205
rect 942 196 944 200
rect 948 196 950 200
rect 942 195 950 196
rect 952 204 959 205
rect 952 200 954 204
rect 958 200 959 204
rect 952 195 959 200
rect 1103 189 1118 190
rect 1107 185 1118 189
rect 1103 184 1118 185
rect 1120 189 1140 190
rect 1120 185 1136 189
rect 1120 184 1140 185
rect 1147 189 1157 190
rect 1147 185 1149 189
rect 1153 185 1157 189
rect 1147 184 1157 185
rect 1159 189 1178 190
rect 1159 185 1166 189
rect 1170 185 1178 189
rect 1159 184 1178 185
rect 1180 189 1188 190
rect 1180 185 1183 189
rect 1187 185 1188 189
rect 1180 184 1188 185
rect 1201 189 1211 190
rect 1201 185 1203 189
rect 1207 185 1211 189
rect 1201 184 1211 185
rect 1213 189 1232 190
rect 1213 185 1220 189
rect 1224 185 1232 189
rect 1213 184 1232 185
rect 1234 189 1242 190
rect 1234 185 1237 189
rect 1241 185 1242 189
rect 1234 184 1242 185
rect 1257 189 1267 190
rect 1257 185 1259 189
rect 1263 185 1267 189
rect 1257 184 1267 185
rect 1269 189 1288 190
rect 1269 185 1276 189
rect 1280 185 1288 189
rect 1269 184 1288 185
rect 1290 189 1298 190
rect 1290 185 1293 189
rect 1297 185 1298 189
rect 1290 184 1298 185
rect 1311 189 1321 190
rect 1311 185 1313 189
rect 1317 185 1321 189
rect 1311 184 1321 185
rect 1323 189 1342 190
rect 1323 185 1330 189
rect 1334 185 1342 189
rect 1323 184 1342 185
rect 1344 189 1352 190
rect 1344 185 1347 189
rect 1351 185 1352 189
rect 1344 184 1352 185
rect 1010 146 1041 147
rect 1010 142 1015 146
rect 1019 142 1041 146
rect 1010 141 1041 142
rect 1043 142 1059 147
rect 1065 142 1078 147
rect 1043 141 1078 142
rect 1098 146 1113 147
rect 1102 142 1113 146
rect 1098 141 1113 142
rect 1115 146 1135 147
rect 1115 142 1131 146
rect 1115 141 1135 142
rect 1142 146 1152 147
rect 1142 142 1144 146
rect 1148 142 1152 146
rect 1142 141 1152 142
rect 1154 146 1173 147
rect 1154 142 1161 146
rect 1165 142 1173 146
rect 1154 141 1173 142
rect 1175 146 1183 147
rect 1175 142 1178 146
rect 1182 142 1183 146
rect 1175 141 1183 142
rect 1196 146 1206 147
rect 1196 142 1198 146
rect 1202 142 1206 146
rect 1196 141 1206 142
rect 1208 146 1227 147
rect 1208 142 1215 146
rect 1219 142 1227 146
rect 1208 141 1227 142
rect 1229 146 1237 147
rect 1229 142 1232 146
rect 1236 142 1237 146
rect 1229 141 1237 142
rect 1252 146 1262 147
rect 1252 142 1254 146
rect 1258 142 1262 146
rect 1252 141 1262 142
rect 1264 146 1283 147
rect 1264 142 1271 146
rect 1275 142 1283 146
rect 1264 141 1283 142
rect 1285 146 1293 147
rect 1285 142 1288 146
rect 1292 142 1293 146
rect 1285 141 1293 142
rect 1306 146 1316 147
rect 1306 142 1308 146
rect 1312 142 1316 146
rect 1306 141 1316 142
rect 1318 146 1337 147
rect 1318 142 1325 146
rect 1329 142 1337 146
rect 1318 141 1337 142
rect 1339 146 1347 147
rect 1339 142 1342 146
rect 1346 142 1347 146
rect 1339 141 1347 142
rect 147 106 155 109
rect 130 101 135 106
rect 128 100 135 101
rect 128 96 129 100
rect 133 96 135 100
rect 128 95 135 96
rect 130 88 135 95
rect 137 88 142 106
rect 144 97 155 106
rect 157 103 162 109
rect 803 111 811 114
rect 476 108 484 111
rect 459 103 464 108
rect 157 102 164 103
rect 157 98 159 102
rect 163 98 164 102
rect 157 97 164 98
rect 457 102 464 103
rect 457 98 458 102
rect 462 98 464 102
rect 457 97 464 98
rect 144 93 153 97
rect 144 89 147 93
rect 151 89 153 93
rect 144 88 153 89
rect 459 90 464 97
rect 466 90 471 108
rect 473 99 484 108
rect 486 105 491 111
rect 786 106 791 111
rect 784 105 791 106
rect 486 104 493 105
rect 486 100 488 104
rect 492 100 493 104
rect 784 101 785 105
rect 789 101 791 105
rect 784 100 791 101
rect 486 99 493 100
rect 473 95 482 99
rect 473 91 476 95
rect 480 91 482 95
rect 786 93 791 100
rect 793 93 798 111
rect 800 102 811 111
rect 813 108 818 114
rect 813 107 820 108
rect 813 103 815 107
rect 819 103 820 107
rect 813 102 820 103
rect 800 98 809 102
rect 800 94 803 98
rect 807 94 809 98
rect 800 93 809 94
rect 473 90 482 91
rect 340 61 346 63
rect 331 56 336 61
rect 329 55 336 56
rect 329 51 330 55
rect 334 51 336 55
rect 329 48 336 51
rect 329 44 330 48
rect 334 44 336 48
rect 329 43 336 44
rect 338 60 346 61
rect 338 56 340 60
rect 344 56 346 60
rect 338 50 346 56
rect 348 62 356 63
rect 348 58 350 62
rect 354 58 356 62
rect 348 55 356 58
rect 348 51 350 55
rect 354 51 356 55
rect 348 50 356 51
rect 358 62 365 63
rect 358 58 360 62
rect 364 58 365 62
rect 433 61 439 63
rect 358 50 365 58
rect 424 56 429 61
rect 422 55 429 56
rect 422 51 423 55
rect 427 51 429 55
rect 338 43 344 50
rect 422 48 429 51
rect 422 44 423 48
rect 427 44 429 48
rect 422 43 429 44
rect 431 60 439 61
rect 431 56 433 60
rect 437 56 439 60
rect 431 50 439 56
rect 441 62 449 63
rect 441 58 443 62
rect 447 58 449 62
rect 441 55 449 58
rect 441 51 443 55
rect 447 51 449 55
rect 441 50 449 51
rect 451 62 458 63
rect 451 58 453 62
rect 457 58 458 62
rect 520 61 526 63
rect 451 50 458 58
rect 511 56 516 61
rect 509 55 516 56
rect 509 51 510 55
rect 514 51 516 55
rect 431 43 437 50
rect 509 48 516 51
rect 509 44 510 48
rect 514 44 516 48
rect 509 43 516 44
rect 518 60 526 61
rect 518 56 520 60
rect 524 56 526 60
rect 518 50 526 56
rect 528 62 536 63
rect 528 58 530 62
rect 534 58 536 62
rect 528 55 536 58
rect 528 51 530 55
rect 534 51 536 55
rect 528 50 536 51
rect 538 62 545 63
rect 538 58 540 62
rect 544 58 545 62
rect 538 50 545 58
rect 518 43 524 50
rect 1102 47 1117 48
rect 1106 43 1117 47
rect 1102 42 1117 43
rect 1119 47 1139 48
rect 1119 43 1135 47
rect 1119 42 1139 43
rect 1146 47 1156 48
rect 1146 43 1148 47
rect 1152 43 1156 47
rect 1146 42 1156 43
rect 1158 47 1177 48
rect 1158 43 1165 47
rect 1169 43 1177 47
rect 1158 42 1177 43
rect 1179 47 1187 48
rect 1179 43 1182 47
rect 1186 43 1187 47
rect 1179 42 1187 43
rect 1200 47 1210 48
rect 1200 43 1202 47
rect 1206 43 1210 47
rect 1200 42 1210 43
rect 1212 47 1231 48
rect 1212 43 1219 47
rect 1223 43 1231 47
rect 1212 42 1231 43
rect 1233 47 1241 48
rect 1233 43 1236 47
rect 1240 43 1241 47
rect 1233 42 1241 43
rect 1256 47 1266 48
rect 1256 43 1258 47
rect 1262 43 1266 47
rect 1256 42 1266 43
rect 1268 47 1287 48
rect 1268 43 1275 47
rect 1279 43 1287 47
rect 1268 42 1287 43
rect 1289 47 1297 48
rect 1289 43 1292 47
rect 1296 43 1297 47
rect 1289 42 1297 43
rect 1310 47 1320 48
rect 1310 43 1312 47
rect 1316 43 1320 47
rect 1310 42 1320 43
rect 1322 47 1341 48
rect 1322 43 1329 47
rect 1333 43 1341 47
rect 1322 42 1341 43
rect 1343 47 1351 48
rect 1343 43 1346 47
rect 1350 43 1351 47
rect 1343 42 1351 43
<< metal1 >>
rect 33 458 474 462
rect 33 436 37 458
rect 516 456 778 460
rect 115 449 116 452
rect 516 454 520 456
rect 467 451 520 454
rect 331 449 457 450
rect 530 449 574 451
rect 115 448 457 449
rect 110 447 457 448
rect 524 448 574 449
rect 623 448 667 451
rect 710 450 754 451
rect 710 448 762 450
rect 524 447 762 448
rect 110 445 536 447
rect 110 441 134 445
rect 138 441 144 445
rect 148 441 221 445
rect 225 441 231 445
rect 235 441 314 445
rect 318 441 324 445
rect 328 444 536 445
rect 328 441 334 444
rect 530 443 536 444
rect 540 443 546 447
rect 550 444 629 447
rect 550 443 574 444
rect 623 443 629 444
rect 633 443 639 447
rect 643 444 716 447
rect 643 443 667 444
rect 710 443 716 444
rect 720 443 726 447
rect 730 444 762 447
rect 730 443 754 444
rect 774 441 778 456
rect 951 452 1366 455
rect 951 451 1002 452
rect 994 441 999 444
rect 114 431 115 435
rect 119 431 134 435
rect 114 424 126 428
rect 121 419 126 424
rect 130 427 134 431
rect 138 433 150 436
rect 138 430 145 433
rect 149 429 150 433
rect 201 431 202 435
rect 206 431 221 435
rect 145 428 150 429
rect 130 423 142 427
rect 138 419 142 423
rect 121 415 128 419
rect 132 415 135 419
rect 114 402 118 411
rect 122 407 127 411
rect 138 404 142 415
rect 146 414 150 428
rect 202 424 213 428
rect 208 419 213 424
rect 217 427 221 431
rect 225 433 237 436
rect 225 430 232 433
rect 236 429 237 433
rect 294 431 295 435
rect 299 431 314 435
rect 232 428 237 429
rect 217 423 229 427
rect 225 419 229 423
rect 208 415 215 419
rect 219 415 222 419
rect 146 411 175 414
rect 146 410 150 411
rect 107 398 118 402
rect 125 402 142 404
rect 129 400 142 402
rect 145 409 150 410
rect 149 405 150 409
rect 145 402 150 405
rect 125 395 129 398
rect 149 398 150 402
rect 145 397 150 398
rect 114 391 115 395
rect 119 391 120 395
rect 114 385 120 391
rect 125 390 129 391
rect 134 393 135 397
rect 139 393 140 397
rect 134 385 140 393
rect 110 381 144 385
rect 148 381 154 385
rect 110 377 154 381
rect 111 370 115 377
rect 171 375 175 411
rect 201 401 205 411
rect 209 407 214 411
rect 225 404 229 415
rect 233 410 237 428
rect 295 424 306 428
rect 301 419 306 424
rect 310 427 314 431
rect 318 433 330 436
rect 534 435 546 438
rect 318 430 325 433
rect 329 429 330 433
rect 343 429 515 433
rect 520 429 521 433
rect 534 431 535 435
rect 539 432 546 435
rect 550 433 565 437
rect 569 433 570 437
rect 627 435 639 438
rect 534 430 539 431
rect 325 428 330 429
rect 310 423 322 427
rect 318 419 322 423
rect 301 415 308 419
rect 312 415 315 419
rect 198 398 205 401
rect 212 402 229 404
rect 216 400 229 402
rect 232 409 237 410
rect 236 405 237 409
rect 232 402 237 405
rect 212 395 216 398
rect 236 400 237 402
rect 236 398 243 400
rect 232 397 243 398
rect 294 401 298 411
rect 302 407 307 411
rect 318 404 322 415
rect 326 410 330 428
rect 534 423 538 430
rect 550 429 554 433
rect 627 431 628 435
rect 632 432 639 435
rect 643 433 658 437
rect 662 433 663 437
rect 714 435 726 438
rect 774 437 980 441
rect 627 430 632 431
rect 478 419 538 423
rect 534 412 538 419
rect 542 425 554 429
rect 558 427 569 430
rect 542 421 546 425
rect 558 421 563 427
rect 549 417 552 421
rect 556 417 563 421
rect 627 419 631 430
rect 643 429 647 433
rect 714 431 715 435
rect 719 432 726 435
rect 730 433 745 437
rect 749 433 750 437
rect 714 430 719 431
rect 534 411 539 412
rect 291 398 298 401
rect 305 402 322 404
rect 309 400 322 402
rect 325 409 330 410
rect 329 405 330 409
rect 343 407 516 410
rect 534 407 535 411
rect 325 402 330 405
rect 201 391 202 395
rect 206 391 207 395
rect 201 385 207 391
rect 212 390 216 391
rect 221 393 222 397
rect 226 393 227 397
rect 305 395 309 398
rect 329 398 330 402
rect 534 404 539 407
rect 534 400 535 404
rect 542 406 546 417
rect 604 416 631 419
rect 557 409 562 413
rect 542 404 559 406
rect 542 402 555 404
rect 534 399 539 400
rect 566 403 570 413
rect 604 404 608 416
rect 566 400 573 403
rect 325 397 330 398
rect 221 385 227 393
rect 294 391 295 395
rect 299 391 300 395
rect 294 385 300 391
rect 305 390 309 391
rect 314 393 315 397
rect 319 393 320 397
rect 544 395 545 399
rect 549 395 550 399
rect 314 385 320 393
rect 343 389 517 392
rect 544 387 550 395
rect 555 397 559 400
rect 627 412 631 416
rect 635 425 647 429
rect 651 429 665 430
rect 651 427 662 429
rect 635 421 639 425
rect 651 421 656 427
rect 642 417 645 421
rect 649 417 656 421
rect 627 411 632 412
rect 627 407 628 411
rect 627 404 632 407
rect 627 400 628 404
rect 635 406 639 417
rect 714 416 718 430
rect 730 429 734 433
rect 650 409 655 413
rect 635 404 652 406
rect 635 402 648 404
rect 627 399 632 400
rect 659 403 663 413
rect 692 412 718 416
rect 722 425 734 429
rect 738 429 752 430
rect 994 429 997 441
rect 1016 433 1019 452
rect 1029 441 1083 444
rect 1061 435 1065 437
rect 738 427 749 429
rect 722 421 726 425
rect 738 421 743 427
rect 753 425 998 429
rect 729 417 732 421
rect 736 417 743 421
rect 1061 418 1065 429
rect 1080 426 1083 441
rect 1099 433 1102 452
rect 1162 433 1165 452
rect 1172 447 1175 452
rect 1216 433 1219 452
rect 1226 447 1229 452
rect 1272 433 1275 452
rect 1282 447 1285 452
rect 1326 433 1329 452
rect 1336 447 1339 452
rect 1080 423 1130 426
rect 659 400 666 403
rect 678 402 679 406
rect 555 392 559 393
rect 564 393 565 397
rect 569 393 570 397
rect 564 387 570 393
rect 637 395 638 399
rect 642 395 643 399
rect 637 387 643 395
rect 648 397 652 400
rect 648 392 652 393
rect 657 393 658 397
rect 662 393 663 397
rect 657 387 663 393
rect 197 381 231 385
rect 235 381 241 385
rect 197 380 241 381
rect 290 381 324 385
rect 328 381 334 385
rect 197 377 224 380
rect 290 377 334 381
rect 530 383 536 387
rect 540 383 574 387
rect 623 383 629 387
rect 633 383 667 387
rect 530 379 574 383
rect 199 370 203 377
rect 236 373 269 376
rect 290 370 294 377
rect 566 375 570 379
rect 585 378 615 381
rect 623 379 667 383
rect 678 382 682 402
rect 524 374 628 375
rect 524 372 650 374
rect 659 372 663 379
rect 692 381 696 412
rect 714 411 719 412
rect 714 407 715 411
rect 702 382 706 402
rect 714 404 719 407
rect 714 400 715 404
rect 722 406 726 417
rect 737 409 742 413
rect 722 404 739 406
rect 722 402 735 404
rect 714 399 719 400
rect 746 404 750 413
rect 1044 414 1047 417
rect 1061 408 1064 418
rect 1116 413 1119 416
rect 746 400 754 404
rect 724 395 725 399
rect 729 395 730 399
rect 724 387 730 395
rect 735 397 739 400
rect 735 392 739 393
rect 744 393 745 397
rect 749 393 750 397
rect 744 387 750 393
rect 710 383 716 387
rect 720 383 754 387
rect 710 379 754 383
rect 748 372 752 379
rect 945 375 949 408
rect 1061 404 1062 408
rect 1061 396 1064 404
rect 1126 403 1130 423
rect 1133 407 1136 429
rect 1146 424 1149 429
rect 1179 424 1182 429
rect 1146 421 1182 424
rect 1148 413 1150 416
rect 1162 414 1166 416
rect 1170 414 1171 416
rect 1162 413 1171 414
rect 1133 403 1134 407
rect 1162 405 1165 413
rect 1179 412 1182 421
rect 1200 424 1203 429
rect 1233 424 1236 429
rect 1200 421 1236 424
rect 1256 424 1259 429
rect 1289 424 1292 429
rect 1256 421 1292 424
rect 1310 424 1313 429
rect 1343 424 1346 429
rect 1310 421 1346 424
rect 1186 412 1189 421
rect 1200 416 1207 417
rect 1200 414 1204 416
rect 1221 412 1225 415
rect 1179 409 1189 412
rect 1162 403 1167 405
rect 1133 395 1136 403
rect 1162 402 1163 403
rect 1179 396 1182 409
rect 1221 408 1224 412
rect 1233 409 1236 421
rect 1289 420 1292 421
rect 1257 413 1260 416
rect 1233 406 1252 409
rect 1233 396 1236 406
rect 1281 410 1284 412
rect 1269 402 1272 408
rect 1283 406 1284 410
rect 1281 405 1284 406
rect 1246 399 1272 402
rect 1289 396 1292 416
rect 1313 412 1314 415
rect 1332 416 1338 417
rect 1332 414 1335 416
rect 1313 403 1316 412
rect 1343 411 1346 421
rect 1315 399 1316 403
rect 1343 396 1346 407
rect 1027 386 1030 392
rect 1099 386 1102 391
rect 1145 386 1148 392
rect 1199 386 1202 392
rect 1255 386 1258 392
rect 1309 386 1312 392
rect 1003 383 1348 386
rect 762 372 964 375
rect 306 371 964 372
rect 306 370 694 371
rect 2 369 229 370
rect 242 369 694 370
rect 2 368 694 369
rect 2 366 367 368
rect 2 362 38 366
rect 42 362 52 366
rect 56 362 66 366
rect 70 363 149 366
rect 70 362 133 363
rect 2 251 6 362
rect 22 361 37 362
rect 36 342 40 349
rect 36 341 41 342
rect 36 337 37 341
rect 44 341 48 362
rect 51 356 64 357
rect 51 352 54 356
rect 58 352 60 356
rect 51 351 64 352
rect 51 344 57 351
rect 67 345 71 362
rect 137 362 149 363
rect 153 363 233 366
rect 153 362 217 363
rect 114 351 126 357
rect 133 356 137 359
rect 221 362 233 363
rect 237 362 270 366
rect 274 362 284 366
rect 288 362 298 366
rect 302 364 367 366
rect 371 364 381 368
rect 385 364 395 368
rect 399 365 478 368
rect 399 364 462 365
rect 302 362 337 364
rect 147 353 169 357
rect 173 353 174 357
rect 198 356 210 357
rect 147 352 151 353
rect 133 351 137 352
rect 114 348 119 351
rect 114 347 115 348
rect 44 337 47 341
rect 51 337 52 341
rect 56 337 57 341
rect 61 337 62 341
rect 67 340 71 341
rect 106 344 115 347
rect 140 348 151 352
rect 198 352 203 356
rect 207 352 210 356
rect 198 351 210 352
rect 217 356 221 359
rect 231 353 253 357
rect 257 353 258 357
rect 231 352 235 353
rect 217 351 221 352
rect 140 344 144 348
rect 158 345 159 349
rect 163 345 174 349
rect 36 336 41 337
rect 36 328 40 336
rect 56 332 62 337
rect 43 328 44 332
rect 48 328 62 332
rect 68 330 72 333
rect 106 330 109 344
rect 114 343 119 344
rect 123 342 144 344
rect 36 319 40 324
rect 36 318 41 319
rect 36 314 37 318
rect 41 314 48 317
rect 36 311 48 314
rect 52 315 56 328
rect 115 338 123 339
rect 127 340 144 342
rect 115 335 127 338
rect 68 324 72 326
rect 59 320 63 324
rect 67 320 72 324
rect 59 319 72 320
rect 115 323 119 335
rect 140 333 144 340
rect 148 338 149 342
rect 153 341 154 342
rect 153 338 165 341
rect 148 337 165 338
rect 161 334 165 337
rect 161 333 166 334
rect 129 327 135 332
rect 140 329 152 333
rect 156 329 157 333
rect 161 329 162 333
rect 129 325 131 327
rect 122 323 131 325
rect 161 328 166 329
rect 170 329 174 345
rect 198 348 203 351
rect 198 344 199 348
rect 224 348 235 352
rect 224 344 228 348
rect 242 345 243 349
rect 247 345 258 349
rect 198 343 203 344
rect 207 342 228 344
rect 199 338 207 339
rect 211 340 228 342
rect 199 335 211 338
rect 161 324 165 328
rect 122 319 135 323
rect 141 320 165 324
rect 170 325 172 329
rect 115 318 119 319
rect 141 318 145 320
rect 52 311 66 315
rect 70 311 71 315
rect 128 311 129 315
rect 133 311 134 315
rect 170 316 174 325
rect 199 323 203 335
rect 224 333 228 340
rect 232 338 233 342
rect 237 341 238 342
rect 237 338 249 341
rect 232 337 249 338
rect 245 334 249 337
rect 245 333 250 334
rect 213 327 219 332
rect 224 329 236 333
rect 240 329 241 333
rect 245 329 246 333
rect 213 325 215 327
rect 206 323 215 325
rect 245 328 250 329
rect 245 324 249 328
rect 206 319 219 323
rect 225 320 249 324
rect 199 318 203 319
rect 225 318 229 320
rect 141 313 145 314
rect 150 312 151 316
rect 155 312 174 316
rect 128 306 134 311
rect 212 311 213 315
rect 217 311 218 315
rect 254 316 258 345
rect 268 342 272 349
rect 268 341 273 342
rect 268 337 269 341
rect 276 341 280 362
rect 283 356 296 357
rect 283 352 286 356
rect 290 352 292 356
rect 283 351 296 352
rect 283 344 289 351
rect 299 345 303 362
rect 276 337 279 341
rect 283 337 284 341
rect 288 337 289 341
rect 293 337 294 341
rect 299 340 303 341
rect 268 336 273 337
rect 268 328 272 336
rect 288 332 294 337
rect 275 328 276 332
rect 280 328 294 332
rect 300 331 304 333
rect 225 313 229 314
rect 234 312 235 316
rect 239 312 258 316
rect 262 325 272 328
rect 262 313 265 325
rect 212 306 218 311
rect 268 319 272 325
rect 268 318 273 319
rect 268 314 269 318
rect 273 314 280 317
rect 268 311 280 314
rect 284 315 288 328
rect 300 324 304 327
rect 291 320 295 324
rect 299 320 304 324
rect 291 319 304 320
rect 284 311 298 315
rect 302 311 303 315
rect 35 302 38 306
rect 42 302 48 306
rect 52 302 116 306
rect 120 302 169 306
rect 173 302 200 306
rect 204 302 253 306
rect 257 302 270 306
rect 274 302 280 306
rect 284 305 308 306
rect 284 302 302 305
rect 21 299 302 302
rect 21 298 308 299
rect 125 296 169 298
rect 125 292 131 296
rect 135 292 159 296
rect 163 292 169 296
rect 129 284 135 292
rect 129 280 130 284
rect 134 280 135 284
rect 140 284 144 285
rect 149 284 155 292
rect 149 280 150 284
rect 154 280 155 284
rect 160 284 165 287
rect 164 280 165 284
rect 140 277 144 280
rect 160 279 165 280
rect 140 273 157 277
rect 129 261 133 271
rect 137 266 142 270
rect 153 269 157 273
rect 137 258 143 262
rect 147 258 150 262
rect 1 231 6 251
rect 137 252 141 258
rect 153 254 157 265
rect 124 249 141 252
rect 145 250 157 254
rect 161 275 322 279
rect 145 246 149 250
rect 161 249 165 275
rect 331 253 335 362
rect 365 344 369 351
rect 365 343 370 344
rect 365 339 366 343
rect 373 343 377 364
rect 380 358 393 359
rect 380 354 383 358
rect 387 354 389 358
rect 380 353 393 354
rect 380 346 386 353
rect 396 347 400 364
rect 466 364 478 365
rect 482 365 562 368
rect 482 364 546 365
rect 443 353 455 359
rect 462 358 466 361
rect 550 364 562 365
rect 566 364 599 368
rect 603 364 613 368
rect 617 364 627 368
rect 631 367 694 368
rect 698 367 708 371
rect 712 367 722 371
rect 726 368 805 371
rect 726 367 789 368
rect 631 364 667 367
rect 476 355 498 359
rect 502 355 503 359
rect 518 358 539 359
rect 476 354 480 355
rect 462 353 466 354
rect 443 350 448 353
rect 443 349 444 350
rect 373 339 376 343
rect 380 339 381 343
rect 385 339 386 343
rect 390 339 391 343
rect 396 342 400 343
rect 435 346 444 349
rect 469 350 480 354
rect 518 354 532 358
rect 536 354 539 358
rect 518 353 539 354
rect 546 358 550 361
rect 560 355 582 359
rect 586 355 587 359
rect 560 354 564 355
rect 546 353 550 354
rect 469 346 473 350
rect 487 347 488 351
rect 492 347 503 351
rect 365 338 370 339
rect 365 330 369 338
rect 385 334 391 339
rect 372 330 373 334
rect 377 330 391 334
rect 397 332 401 335
rect 435 332 438 346
rect 443 345 448 346
rect 452 344 473 346
rect 365 321 369 326
rect 365 320 370 321
rect 365 316 366 320
rect 370 316 377 319
rect 365 313 377 316
rect 381 317 385 330
rect 444 340 452 341
rect 456 342 473 344
rect 444 337 456 340
rect 397 326 401 328
rect 388 322 392 326
rect 396 322 401 326
rect 388 321 401 322
rect 444 325 448 337
rect 469 335 473 342
rect 477 340 478 344
rect 482 343 483 344
rect 482 340 494 343
rect 477 339 494 340
rect 490 336 494 339
rect 490 335 495 336
rect 458 329 464 334
rect 469 331 481 335
rect 485 331 486 335
rect 490 331 491 335
rect 458 327 460 329
rect 451 325 460 327
rect 490 330 495 331
rect 499 331 503 347
rect 527 350 532 353
rect 527 346 528 350
rect 553 350 564 354
rect 553 346 557 350
rect 571 347 572 351
rect 576 347 589 351
rect 527 345 532 346
rect 536 344 557 346
rect 528 340 536 341
rect 540 342 557 344
rect 528 337 540 340
rect 490 326 494 330
rect 451 321 464 325
rect 470 322 494 326
rect 499 327 501 331
rect 444 320 448 321
rect 470 320 474 322
rect 381 313 395 317
rect 399 313 400 317
rect 457 313 458 317
rect 462 313 463 317
rect 499 318 503 327
rect 528 325 532 337
rect 553 335 557 342
rect 561 340 562 344
rect 566 343 567 344
rect 566 340 578 343
rect 561 339 578 340
rect 574 336 578 339
rect 574 335 579 336
rect 542 329 548 334
rect 553 331 565 335
rect 569 331 570 335
rect 574 331 575 335
rect 542 327 544 329
rect 535 325 544 327
rect 574 330 579 331
rect 574 326 578 330
rect 535 321 548 325
rect 554 322 578 326
rect 528 320 532 321
rect 554 320 558 322
rect 470 315 474 316
rect 479 314 480 318
rect 484 314 503 318
rect 457 308 463 313
rect 541 313 542 317
rect 546 313 547 317
rect 583 318 587 347
rect 597 344 601 351
rect 597 343 602 344
rect 597 339 598 343
rect 605 343 609 364
rect 612 358 625 359
rect 612 354 615 358
rect 619 354 621 358
rect 612 353 625 354
rect 612 346 618 353
rect 628 347 632 364
rect 605 339 608 343
rect 612 339 613 343
rect 617 339 618 343
rect 622 339 623 343
rect 628 342 632 343
rect 597 338 602 339
rect 597 330 601 338
rect 617 334 623 339
rect 604 330 605 334
rect 609 330 623 334
rect 629 333 633 335
rect 554 315 558 316
rect 563 314 564 318
rect 568 314 587 318
rect 591 327 601 330
rect 591 315 594 327
rect 541 308 547 313
rect 597 321 601 327
rect 597 320 602 321
rect 597 316 598 320
rect 602 316 609 319
rect 597 313 609 316
rect 613 317 617 330
rect 629 326 633 329
rect 620 322 624 326
rect 628 322 633 326
rect 620 321 633 322
rect 613 313 627 317
rect 631 313 632 317
rect 364 304 367 308
rect 371 304 377 308
rect 381 304 445 308
rect 449 304 498 308
rect 502 304 529 308
rect 533 304 582 308
rect 586 304 599 308
rect 603 304 609 308
rect 613 307 637 308
rect 613 304 629 307
rect 364 303 629 304
rect 349 301 629 303
rect 635 301 637 307
rect 349 300 637 301
rect 349 299 365 300
rect 454 298 498 300
rect 454 294 460 298
rect 464 294 488 298
rect 492 294 498 298
rect 458 286 464 294
rect 458 282 459 286
rect 463 282 464 286
rect 469 286 473 287
rect 478 286 484 294
rect 478 282 479 286
rect 483 282 484 286
rect 489 286 494 289
rect 493 282 494 286
rect 469 279 473 282
rect 489 281 494 282
rect 351 275 419 279
rect 469 275 486 279
rect 458 263 462 273
rect 466 268 471 272
rect 482 271 486 275
rect 466 260 472 264
rect 476 260 479 264
rect 160 248 165 249
rect 129 242 130 246
rect 134 242 149 246
rect 152 244 160 246
rect 164 244 165 248
rect 152 242 165 244
rect 147 236 148 239
rect 125 235 148 236
rect 152 236 153 239
rect 152 235 159 236
rect 125 232 159 235
rect 163 232 169 236
rect 125 231 169 232
rect 330 233 335 253
rect 466 254 470 260
rect 482 256 486 267
rect 453 251 470 254
rect 474 252 486 256
rect 490 275 494 281
rect 490 272 641 275
rect 645 272 646 275
rect 474 248 478 252
rect 490 251 494 272
rect 658 256 662 364
rect 692 347 696 354
rect 692 346 697 347
rect 692 342 693 346
rect 700 346 704 367
rect 707 361 720 362
rect 707 357 710 361
rect 714 357 716 361
rect 707 356 720 357
rect 707 349 713 356
rect 723 350 727 367
rect 793 367 805 368
rect 809 368 889 371
rect 809 367 873 368
rect 770 356 782 362
rect 789 361 793 364
rect 877 367 889 368
rect 893 367 926 371
rect 930 367 940 371
rect 944 367 954 371
rect 958 367 964 371
rect 803 358 825 362
rect 829 358 830 362
rect 843 361 866 362
rect 803 357 807 358
rect 843 357 859 361
rect 863 357 866 361
rect 789 356 793 357
rect 770 353 775 356
rect 770 352 771 353
rect 700 342 703 346
rect 707 342 708 346
rect 712 342 713 346
rect 717 342 718 346
rect 723 345 727 346
rect 692 341 697 342
rect 692 333 696 341
rect 712 337 718 342
rect 699 333 700 337
rect 704 333 718 337
rect 724 335 728 338
rect 692 324 696 329
rect 692 323 697 324
rect 692 319 693 323
rect 697 319 704 322
rect 692 316 704 319
rect 708 320 712 333
rect 724 329 728 331
rect 715 325 719 329
rect 723 325 728 329
rect 715 324 728 325
rect 708 316 722 320
rect 726 316 727 320
rect 751 318 755 347
rect 762 349 771 352
rect 796 353 807 357
rect 796 349 800 353
rect 814 350 815 354
rect 819 350 830 354
rect 762 335 765 349
rect 770 348 775 349
rect 779 347 800 349
rect 771 343 779 344
rect 783 345 800 347
rect 771 340 783 343
rect 771 328 775 340
rect 796 338 800 345
rect 804 343 805 347
rect 809 346 810 347
rect 809 343 821 346
rect 804 342 821 343
rect 817 339 821 342
rect 817 338 822 339
rect 785 332 791 337
rect 796 334 808 338
rect 812 334 813 338
rect 817 334 818 338
rect 785 330 787 332
rect 778 328 787 330
rect 817 333 822 334
rect 826 334 830 350
rect 817 329 821 333
rect 778 324 791 328
rect 797 325 821 329
rect 826 330 828 334
rect 771 323 775 324
rect 797 323 801 325
rect 751 314 752 318
rect 784 316 785 320
rect 789 316 790 320
rect 826 321 830 330
rect 797 318 801 319
rect 806 317 807 321
rect 811 317 830 321
rect 837 318 840 349
rect 784 311 790 316
rect 844 311 848 357
rect 854 356 866 357
rect 873 361 877 364
rect 887 358 909 362
rect 913 358 914 362
rect 887 357 891 358
rect 873 356 877 357
rect 854 353 859 356
rect 854 349 855 353
rect 880 353 891 357
rect 880 349 884 353
rect 898 350 899 354
rect 903 350 914 354
rect 854 348 859 349
rect 863 347 884 349
rect 855 343 863 344
rect 867 345 884 347
rect 855 340 867 343
rect 855 328 859 340
rect 880 338 884 345
rect 888 343 889 347
rect 893 346 894 347
rect 893 343 905 346
rect 888 342 905 343
rect 901 339 905 342
rect 901 338 906 339
rect 869 332 875 337
rect 880 334 892 338
rect 896 334 897 338
rect 901 334 902 338
rect 869 330 871 332
rect 862 328 871 330
rect 901 333 906 334
rect 901 329 905 333
rect 862 324 875 328
rect 881 325 905 329
rect 855 323 859 324
rect 881 323 885 325
rect 868 316 869 320
rect 873 316 874 320
rect 910 321 914 350
rect 924 347 928 354
rect 924 346 929 347
rect 924 342 925 346
rect 932 346 936 367
rect 939 361 952 362
rect 939 357 942 361
rect 946 357 948 361
rect 939 356 952 357
rect 939 349 945 356
rect 955 350 959 367
rect 932 342 935 346
rect 939 342 940 346
rect 944 342 945 346
rect 949 342 950 346
rect 955 345 959 346
rect 924 341 929 342
rect 924 333 928 341
rect 944 337 950 342
rect 931 333 932 337
rect 936 333 950 337
rect 956 336 960 338
rect 881 318 885 319
rect 890 317 891 321
rect 895 317 914 321
rect 918 330 928 333
rect 918 318 921 330
rect 868 311 874 316
rect 924 324 928 330
rect 924 323 929 324
rect 924 319 925 323
rect 929 319 936 322
rect 924 316 936 319
rect 940 320 944 333
rect 956 329 960 332
rect 1003 330 1007 383
rect 1171 380 1176 383
rect 1277 380 1281 383
rect 1103 377 1352 380
rect 1103 372 1106 377
rect 1149 371 1152 377
rect 1203 371 1206 377
rect 1259 371 1262 377
rect 1313 371 1316 377
rect 1137 360 1140 368
rect 1137 356 1138 360
rect 947 325 951 329
rect 955 325 960 329
rect 947 324 960 325
rect 971 326 1007 330
rect 940 316 954 320
rect 958 316 959 320
rect 691 310 694 311
rect 689 307 694 310
rect 698 307 704 311
rect 708 307 772 311
rect 776 307 825 311
rect 829 307 856 311
rect 860 307 909 311
rect 913 307 926 311
rect 930 307 936 311
rect 940 307 964 311
rect 971 307 975 326
rect 689 305 975 307
rect 676 303 975 305
rect 676 302 693 303
rect 676 301 692 302
rect 781 301 825 303
rect 781 297 787 301
rect 791 297 815 301
rect 819 297 825 301
rect 785 289 791 297
rect 785 285 786 289
rect 790 285 791 289
rect 796 289 800 290
rect 805 289 811 297
rect 805 285 806 289
rect 810 285 811 289
rect 816 289 821 292
rect 820 285 821 289
rect 677 272 744 275
rect 748 272 749 275
rect 489 250 494 251
rect 458 244 459 248
rect 463 244 478 248
rect 481 246 489 248
rect 493 246 494 250
rect 481 244 494 246
rect 476 238 477 241
rect 454 237 477 238
rect 481 238 482 241
rect 481 237 488 238
rect 454 234 488 237
rect 492 234 498 238
rect 454 233 498 234
rect 1 228 169 231
rect 1 227 129 228
rect 307 227 322 231
rect 126 224 129 227
rect 330 230 498 233
rect 657 236 662 256
rect 754 244 758 284
rect 796 282 800 285
rect 816 284 821 285
rect 796 278 813 282
rect 766 250 769 277
rect 785 266 789 276
rect 793 271 798 275
rect 809 274 813 278
rect 793 263 799 267
rect 803 263 806 267
rect 793 257 797 263
rect 809 259 813 270
rect 780 254 797 257
rect 801 255 813 259
rect 817 280 821 284
rect 817 277 829 280
rect 801 251 805 255
rect 817 254 821 277
rect 837 256 840 271
rect 816 253 821 254
rect 785 247 786 251
rect 790 247 805 251
rect 808 249 816 251
rect 820 249 821 253
rect 808 247 821 249
rect 803 241 804 244
rect 754 239 758 240
rect 781 240 804 241
rect 808 241 809 244
rect 836 243 841 256
rect 808 240 815 241
rect 781 237 815 240
rect 819 237 825 241
rect 781 236 825 237
rect 987 241 990 326
rect 1086 322 1090 350
rect 1120 347 1123 350
rect 1137 334 1140 356
rect 1183 354 1186 367
rect 1183 351 1193 354
rect 1225 351 1228 355
rect 1237 357 1240 367
rect 1237 354 1256 357
rect 1285 357 1288 358
rect 1152 347 1154 350
rect 1174 347 1175 350
rect 1183 342 1186 351
rect 1150 339 1186 342
rect 1150 334 1153 339
rect 1183 334 1186 339
rect 1190 342 1193 351
rect 1204 347 1208 349
rect 1225 348 1229 351
rect 1204 346 1211 347
rect 1237 342 1240 354
rect 1287 353 1288 357
rect 1285 351 1288 353
rect 1261 347 1264 350
rect 1293 347 1296 367
rect 1319 360 1320 364
rect 1317 351 1320 360
rect 1347 356 1350 367
rect 1317 348 1318 351
rect 1336 347 1339 349
rect 1336 346 1342 347
rect 1293 342 1296 343
rect 1347 342 1350 352
rect 1204 339 1240 342
rect 1204 334 1207 339
rect 1237 334 1240 339
rect 1260 339 1296 342
rect 1260 334 1263 339
rect 1293 334 1296 339
rect 1314 339 1350 342
rect 1314 334 1317 339
rect 1347 334 1350 339
rect 1089 320 1090 322
rect 1103 311 1106 330
rect 1166 311 1169 330
rect 1176 311 1179 316
rect 1220 311 1223 330
rect 1230 311 1233 316
rect 1276 311 1279 330
rect 1286 311 1289 316
rect 1330 311 1333 330
rect 1340 311 1343 316
rect 1361 311 1366 452
rect 1101 310 1366 311
rect 1000 307 1366 310
rect 1016 288 1019 307
rect 1061 290 1065 292
rect 1099 288 1102 307
rect 1112 299 1142 302
rect 1061 273 1065 284
rect 1044 269 1047 272
rect 1061 263 1064 273
rect 1116 268 1119 271
rect 1061 259 1062 263
rect 1133 262 1136 284
rect 1139 272 1142 299
rect 1162 288 1165 307
rect 1172 302 1175 307
rect 1216 288 1219 307
rect 1226 302 1229 307
rect 1272 288 1275 307
rect 1282 302 1285 307
rect 1326 288 1329 307
rect 1336 302 1339 307
rect 1146 279 1149 284
rect 1179 279 1182 284
rect 1146 276 1182 279
rect 1139 269 1144 272
rect 1148 268 1150 271
rect 1170 268 1171 271
rect 1179 267 1182 276
rect 1200 279 1203 284
rect 1233 279 1236 284
rect 1200 276 1236 279
rect 1256 279 1259 284
rect 1289 279 1292 284
rect 1256 276 1292 279
rect 1310 279 1313 284
rect 1343 279 1346 284
rect 1310 276 1346 279
rect 1186 267 1189 276
rect 1200 271 1207 272
rect 1200 269 1204 271
rect 1221 267 1225 270
rect 1179 264 1189 267
rect 1061 251 1064 259
rect 1133 258 1134 262
rect 1133 250 1136 258
rect 1179 251 1182 264
rect 1221 263 1224 267
rect 1233 264 1236 276
rect 1289 275 1292 276
rect 1257 268 1260 271
rect 1233 261 1252 264
rect 1233 251 1236 261
rect 1281 265 1284 267
rect 1269 257 1272 263
rect 1283 261 1284 265
rect 1281 260 1284 261
rect 1246 254 1272 257
rect 1289 251 1292 271
rect 1313 267 1314 270
rect 1332 271 1338 272
rect 1332 269 1335 271
rect 1313 258 1316 267
rect 1343 266 1346 276
rect 1315 254 1316 258
rect 1343 251 1346 262
rect 1027 241 1030 247
rect 1099 241 1102 246
rect 1145 241 1148 247
rect 1199 241 1202 247
rect 1255 241 1258 247
rect 1309 241 1312 247
rect 987 238 1348 241
rect 657 233 825 236
rect 657 232 781 233
rect 330 229 456 230
rect 786 229 789 233
rect 453 226 456 229
rect 1 220 307 224
rect 1 216 37 220
rect 41 216 51 220
rect 55 216 65 220
rect 69 217 148 220
rect 69 216 132 217
rect 1 105 5 216
rect 35 196 39 203
rect 35 195 40 196
rect 35 191 36 195
rect 43 195 47 216
rect 50 210 63 211
rect 50 206 53 210
rect 57 206 59 210
rect 50 205 63 206
rect 50 198 56 205
rect 66 199 70 216
rect 136 216 148 217
rect 152 217 232 220
rect 152 216 216 217
rect 113 205 125 211
rect 132 210 136 213
rect 220 216 232 217
rect 236 216 269 220
rect 273 216 283 220
rect 287 216 297 220
rect 301 216 307 220
rect 330 222 636 226
rect 330 218 366 222
rect 370 218 380 222
rect 384 218 394 222
rect 398 219 477 222
rect 398 218 461 219
rect 146 207 168 211
rect 172 207 173 211
rect 197 210 209 211
rect 185 207 202 210
rect 146 206 150 207
rect 132 205 136 206
rect 113 202 118 205
rect 113 201 114 202
rect 43 191 46 195
rect 50 191 51 195
rect 55 191 56 195
rect 60 191 61 195
rect 66 194 70 195
rect 105 198 114 201
rect 139 202 150 206
rect 139 198 143 202
rect 157 199 158 203
rect 162 199 173 203
rect 35 190 40 191
rect 35 182 39 190
rect 55 186 61 191
rect 42 182 43 186
rect 47 182 61 186
rect 67 184 71 187
rect 105 184 108 198
rect 113 197 118 198
rect 122 196 143 198
rect 35 173 39 178
rect 35 172 40 173
rect 35 168 36 172
rect 40 168 47 171
rect 35 165 47 168
rect 51 169 55 182
rect 114 192 122 193
rect 126 194 143 196
rect 114 189 126 192
rect 67 178 71 180
rect 58 174 62 178
rect 66 174 71 178
rect 58 173 71 174
rect 114 177 118 189
rect 139 187 143 194
rect 147 192 148 196
rect 152 195 153 196
rect 152 192 164 195
rect 147 191 164 192
rect 160 188 164 191
rect 160 187 165 188
rect 128 181 134 186
rect 139 183 151 187
rect 155 183 156 187
rect 160 183 161 187
rect 128 179 130 181
rect 121 177 130 179
rect 160 182 165 183
rect 169 183 173 199
rect 160 178 164 182
rect 121 173 134 177
rect 140 174 164 178
rect 169 179 171 183
rect 114 172 118 173
rect 140 172 144 174
rect 51 165 65 169
rect 69 165 70 169
rect 127 165 128 169
rect 132 165 133 169
rect 169 170 173 179
rect 140 167 144 168
rect 149 166 150 170
rect 154 166 173 170
rect 185 167 188 207
rect 197 206 202 207
rect 206 206 209 210
rect 197 205 209 206
rect 216 210 220 213
rect 230 207 252 211
rect 256 207 257 211
rect 230 206 234 207
rect 216 205 220 206
rect 197 202 202 205
rect 197 198 198 202
rect 223 202 234 206
rect 223 198 227 202
rect 241 199 242 203
rect 246 199 257 203
rect 197 197 202 198
rect 206 196 227 198
rect 198 192 206 193
rect 210 194 227 196
rect 198 189 210 192
rect 198 177 202 189
rect 223 187 227 194
rect 231 192 232 196
rect 236 195 237 196
rect 236 192 248 195
rect 231 191 248 192
rect 244 188 248 191
rect 244 187 249 188
rect 212 181 218 186
rect 223 183 235 187
rect 239 183 240 187
rect 244 183 245 187
rect 212 179 214 181
rect 205 177 214 179
rect 244 182 249 183
rect 244 178 248 182
rect 205 173 218 177
rect 224 174 248 178
rect 198 172 202 173
rect 224 172 228 174
rect 127 160 133 165
rect 211 165 212 169
rect 216 165 217 169
rect 253 170 257 199
rect 267 196 271 203
rect 267 195 272 196
rect 267 191 268 195
rect 275 195 279 216
rect 282 210 295 211
rect 282 206 285 210
rect 289 206 291 210
rect 282 205 295 206
rect 282 198 288 205
rect 298 199 302 216
rect 275 191 278 195
rect 282 191 283 195
rect 287 191 288 195
rect 292 191 293 195
rect 298 194 302 195
rect 267 190 272 191
rect 267 182 271 190
rect 287 186 293 191
rect 274 182 275 186
rect 279 182 293 186
rect 299 185 303 187
rect 224 167 228 168
rect 233 166 234 170
rect 238 166 257 170
rect 261 179 271 182
rect 261 167 264 179
rect 211 160 217 165
rect 267 173 271 179
rect 267 172 272 173
rect 267 168 268 172
rect 272 168 279 171
rect 267 165 279 168
rect 283 169 287 182
rect 299 178 303 181
rect 290 174 294 178
rect 298 174 303 178
rect 290 173 303 174
rect 283 165 297 169
rect 301 165 302 169
rect 34 156 37 160
rect 41 156 47 160
rect 51 156 115 160
rect 119 156 168 160
rect 172 156 199 160
rect 203 156 252 160
rect 256 156 269 160
rect 273 156 279 160
rect 283 156 302 160
rect 34 153 302 156
rect 34 152 307 153
rect 124 150 168 152
rect 124 146 130 150
rect 134 146 158 150
rect 162 146 168 150
rect 128 138 134 146
rect 128 134 129 138
rect 133 134 134 138
rect 139 138 143 139
rect 148 138 154 146
rect 255 143 296 146
rect 148 134 149 138
rect 153 134 154 138
rect 159 138 164 141
rect 163 134 164 138
rect 139 131 143 134
rect 159 133 164 134
rect 139 127 156 131
rect 128 115 132 125
rect 136 120 141 124
rect 152 123 156 127
rect 136 112 142 116
rect 146 112 149 116
rect 0 85 5 105
rect 136 106 140 112
rect 152 108 156 119
rect 123 103 140 106
rect 144 104 156 108
rect 144 100 148 104
rect 160 103 164 133
rect 252 125 275 128
rect 280 125 281 128
rect 159 102 164 103
rect 128 96 129 100
rect 133 96 148 100
rect 151 98 159 100
rect 163 98 164 102
rect 151 96 164 98
rect 146 90 147 93
rect 124 89 147 90
rect 151 90 152 93
rect 151 89 158 90
rect 124 86 158 89
rect 162 86 168 90
rect 124 85 168 86
rect 0 82 168 85
rect 0 81 124 82
rect 293 42 296 143
rect 305 124 321 128
rect 330 107 334 218
rect 364 198 368 205
rect 364 197 369 198
rect 364 193 365 197
rect 372 197 376 218
rect 379 212 392 213
rect 379 208 382 212
rect 386 208 388 212
rect 379 207 392 208
rect 379 200 385 207
rect 395 201 399 218
rect 465 218 477 219
rect 481 219 561 222
rect 481 218 545 219
rect 442 207 454 213
rect 461 212 465 215
rect 549 218 561 219
rect 565 218 598 222
rect 602 218 612 222
rect 616 218 626 222
rect 630 218 636 222
rect 657 225 963 229
rect 657 221 693 225
rect 697 221 707 225
rect 711 221 721 225
rect 725 222 804 225
rect 725 221 788 222
rect 475 209 497 213
rect 501 209 502 213
rect 526 212 538 213
rect 475 208 479 209
rect 461 207 465 208
rect 442 204 447 207
rect 442 203 443 204
rect 372 193 375 197
rect 379 193 380 197
rect 384 193 385 197
rect 389 193 390 197
rect 395 196 399 197
rect 434 200 443 203
rect 468 204 479 208
rect 526 208 531 212
rect 535 208 538 212
rect 526 207 538 208
rect 545 212 549 215
rect 559 209 581 213
rect 585 209 586 213
rect 559 208 563 209
rect 545 207 549 208
rect 468 200 472 204
rect 486 201 487 205
rect 491 201 502 205
rect 364 192 369 193
rect 364 184 368 192
rect 384 188 390 193
rect 371 184 372 188
rect 376 184 390 188
rect 396 186 400 189
rect 364 175 368 180
rect 364 174 369 175
rect 364 170 365 174
rect 369 170 376 173
rect 364 167 376 170
rect 380 171 384 184
rect 396 180 400 182
rect 387 176 391 180
rect 395 176 400 180
rect 387 175 400 176
rect 380 167 394 171
rect 398 167 399 171
rect 424 169 427 189
rect 434 186 437 200
rect 442 199 447 200
rect 451 198 472 200
rect 443 194 451 195
rect 455 196 472 198
rect 443 191 455 194
rect 443 179 447 191
rect 468 189 472 196
rect 476 194 477 198
rect 481 197 482 198
rect 481 194 493 197
rect 476 193 493 194
rect 489 190 493 193
rect 489 189 494 190
rect 457 183 463 188
rect 468 185 480 189
rect 484 185 485 189
rect 489 185 490 189
rect 457 181 459 183
rect 450 179 459 181
rect 489 184 494 185
rect 498 185 502 201
rect 526 204 531 207
rect 526 200 527 204
rect 552 204 563 208
rect 552 200 556 204
rect 570 201 571 205
rect 575 201 586 205
rect 526 199 531 200
rect 535 198 556 200
rect 527 194 535 195
rect 539 196 556 198
rect 527 191 539 194
rect 489 180 493 184
rect 450 175 463 179
rect 469 176 493 180
rect 498 181 500 185
rect 443 174 447 175
rect 469 174 473 176
rect 456 167 457 171
rect 461 167 462 171
rect 498 172 502 181
rect 527 179 531 191
rect 552 189 556 196
rect 560 194 561 198
rect 565 197 566 198
rect 565 194 577 197
rect 560 193 577 194
rect 573 190 577 193
rect 573 189 578 190
rect 541 183 547 188
rect 552 185 564 189
rect 568 185 569 189
rect 573 185 574 189
rect 541 181 543 183
rect 534 179 543 181
rect 573 184 578 185
rect 573 180 577 184
rect 534 175 547 179
rect 553 176 577 180
rect 527 174 531 175
rect 553 174 557 176
rect 469 169 473 170
rect 478 168 479 172
rect 483 168 502 172
rect 456 162 462 167
rect 540 167 541 171
rect 545 167 546 171
rect 582 172 586 201
rect 596 198 600 205
rect 596 197 601 198
rect 596 193 597 197
rect 604 197 608 218
rect 611 212 624 213
rect 611 208 614 212
rect 618 208 620 212
rect 611 207 624 208
rect 611 200 617 207
rect 627 201 631 218
rect 604 193 607 197
rect 611 193 612 197
rect 616 193 617 197
rect 621 193 622 197
rect 627 196 631 197
rect 596 192 601 193
rect 596 184 600 192
rect 616 188 622 193
rect 603 184 604 188
rect 608 184 622 188
rect 628 187 632 189
rect 553 169 557 170
rect 562 168 563 172
rect 567 168 586 172
rect 590 181 600 184
rect 590 169 593 181
rect 540 162 546 167
rect 596 175 600 181
rect 596 174 601 175
rect 596 170 597 174
rect 601 170 608 173
rect 596 167 608 170
rect 612 171 616 184
rect 628 180 632 183
rect 619 176 623 180
rect 627 176 632 180
rect 619 175 632 176
rect 612 167 626 171
rect 630 167 631 171
rect 363 158 366 162
rect 370 158 376 162
rect 380 158 444 162
rect 448 158 497 162
rect 501 158 528 162
rect 532 158 581 162
rect 585 158 598 162
rect 602 158 608 162
rect 612 158 636 162
rect 344 155 629 158
rect 363 154 629 155
rect 633 154 636 158
rect 453 152 497 154
rect 453 148 459 152
rect 463 148 487 152
rect 491 148 497 152
rect 424 143 427 145
rect 457 140 463 148
rect 424 125 427 139
rect 457 136 458 140
rect 462 136 463 140
rect 468 140 472 141
rect 477 140 483 148
rect 477 136 478 140
rect 482 136 483 140
rect 488 140 493 143
rect 492 136 493 140
rect 468 133 472 136
rect 488 135 493 136
rect 468 129 485 133
rect 329 87 334 107
rect 396 121 424 124
rect 396 95 400 121
rect 457 117 461 127
rect 465 122 470 126
rect 481 125 485 129
rect 465 114 471 118
rect 475 114 478 118
rect 465 108 469 114
rect 481 110 485 121
rect 452 105 469 108
rect 473 106 485 110
rect 473 102 477 106
rect 489 105 493 135
rect 520 131 602 136
rect 657 110 661 221
rect 691 201 695 208
rect 691 200 696 201
rect 691 196 692 200
rect 699 200 703 221
rect 706 215 719 216
rect 706 211 709 215
rect 713 211 715 215
rect 706 210 719 211
rect 706 203 712 210
rect 722 204 726 221
rect 792 221 804 222
rect 808 222 888 225
rect 808 221 872 222
rect 769 210 781 216
rect 788 215 792 218
rect 876 221 888 222
rect 892 221 925 225
rect 929 221 939 225
rect 943 221 953 225
rect 957 221 963 225
rect 802 212 824 216
rect 828 212 829 216
rect 853 215 865 216
rect 802 211 806 212
rect 788 210 792 211
rect 769 207 774 210
rect 769 206 770 207
rect 699 196 702 200
rect 706 196 707 200
rect 711 196 712 200
rect 716 196 717 200
rect 722 199 726 200
rect 761 203 770 206
rect 795 207 806 211
rect 853 211 858 215
rect 862 211 865 215
rect 853 210 865 211
rect 872 215 876 218
rect 886 212 908 216
rect 912 212 913 216
rect 886 211 890 212
rect 872 210 876 211
rect 795 203 799 207
rect 813 204 814 208
rect 818 204 829 208
rect 691 195 696 196
rect 691 187 695 195
rect 711 191 717 196
rect 698 187 699 191
rect 703 187 717 191
rect 723 189 727 192
rect 761 189 764 203
rect 769 202 774 203
rect 778 201 799 203
rect 691 178 695 183
rect 691 177 696 178
rect 691 173 692 177
rect 696 173 703 176
rect 691 170 703 173
rect 707 174 711 187
rect 770 197 778 198
rect 782 199 799 201
rect 770 194 782 197
rect 723 183 727 185
rect 714 179 718 183
rect 722 179 727 183
rect 714 178 727 179
rect 770 182 774 194
rect 795 192 799 199
rect 803 197 804 201
rect 808 200 809 201
rect 808 197 820 200
rect 803 196 820 197
rect 816 193 820 196
rect 816 192 821 193
rect 784 186 790 191
rect 795 188 807 192
rect 811 188 812 192
rect 816 188 817 192
rect 784 184 786 186
rect 770 177 774 178
rect 777 182 786 184
rect 816 187 821 188
rect 825 188 829 204
rect 853 207 858 210
rect 853 203 854 207
rect 879 207 890 211
rect 879 203 883 207
rect 897 204 898 208
rect 902 204 913 208
rect 853 202 858 203
rect 862 201 883 203
rect 854 197 862 198
rect 866 199 883 201
rect 854 194 866 197
rect 816 183 820 187
rect 777 178 790 182
rect 796 179 820 183
rect 825 184 827 188
rect 707 170 721 174
rect 725 170 726 174
rect 777 173 780 178
rect 796 177 800 179
rect 766 169 780 173
rect 783 170 784 174
rect 788 170 789 174
rect 825 175 829 184
rect 854 182 858 194
rect 879 192 883 199
rect 887 197 888 201
rect 892 200 893 201
rect 892 197 904 200
rect 887 196 904 197
rect 900 193 904 196
rect 900 192 905 193
rect 868 186 874 191
rect 879 188 891 192
rect 895 188 896 192
rect 900 188 901 192
rect 868 184 870 186
rect 861 182 870 184
rect 900 187 905 188
rect 900 183 904 187
rect 861 178 874 182
rect 880 179 904 183
rect 854 177 858 178
rect 880 177 884 179
rect 796 172 800 173
rect 805 171 806 175
rect 810 171 829 175
rect 766 165 770 169
rect 783 165 789 170
rect 867 170 868 174
rect 872 170 873 174
rect 909 175 913 204
rect 923 201 927 208
rect 923 200 928 201
rect 923 196 924 200
rect 931 200 935 221
rect 938 215 951 216
rect 938 211 941 215
rect 945 211 947 215
rect 938 210 951 211
rect 938 203 944 210
rect 954 204 958 221
rect 931 196 934 200
rect 938 196 939 200
rect 943 196 944 200
rect 948 196 949 200
rect 954 199 958 200
rect 923 195 928 196
rect 923 187 927 195
rect 943 191 949 196
rect 930 187 931 191
rect 935 187 949 191
rect 955 190 959 192
rect 880 172 884 173
rect 889 171 890 175
rect 894 171 913 175
rect 917 184 927 187
rect 917 172 920 184
rect 867 165 873 170
rect 923 178 927 184
rect 923 177 928 178
rect 923 173 924 177
rect 928 173 935 176
rect 923 170 935 173
rect 939 174 943 187
rect 955 183 959 186
rect 946 179 950 183
rect 954 179 959 183
rect 946 178 959 179
rect 939 170 953 174
rect 957 170 958 174
rect 690 162 693 165
rect 689 161 693 162
rect 697 161 703 165
rect 707 161 771 165
rect 775 161 824 165
rect 828 161 855 165
rect 859 161 908 165
rect 912 161 925 165
rect 929 161 935 165
rect 939 161 963 165
rect 689 159 963 161
rect 670 158 963 159
rect 673 157 963 158
rect 673 156 692 157
rect 780 155 824 157
rect 780 151 786 155
rect 790 151 814 155
rect 818 151 824 155
rect 727 149 731 150
rect 671 131 700 136
rect 488 104 493 105
rect 457 98 458 102
rect 462 98 477 102
rect 480 100 488 102
rect 492 102 493 104
rect 492 100 497 102
rect 480 98 497 100
rect 475 92 476 95
rect 453 91 476 92
rect 480 92 481 95
rect 480 91 487 92
rect 453 88 487 91
rect 491 88 497 92
rect 453 87 497 88
rect 329 84 497 87
rect 656 90 661 110
rect 727 108 731 145
rect 784 143 790 151
rect 784 139 785 143
rect 789 139 790 143
rect 795 143 799 144
rect 804 143 810 151
rect 804 139 805 143
rect 809 139 810 143
rect 815 143 820 146
rect 819 139 820 143
rect 795 136 799 139
rect 815 138 820 139
rect 795 132 812 136
rect 784 120 788 130
rect 792 125 797 129
rect 808 128 812 132
rect 792 117 798 121
rect 802 117 805 121
rect 792 111 796 117
rect 808 113 812 124
rect 779 108 796 111
rect 800 109 812 113
rect 816 133 832 138
rect 800 105 804 109
rect 816 108 820 133
rect 815 107 820 108
rect 784 101 785 105
rect 789 101 804 105
rect 807 103 815 105
rect 819 103 820 107
rect 807 101 820 103
rect 987 99 990 238
rect 1171 235 1176 238
rect 1277 235 1281 238
rect 1103 232 1352 235
rect 1103 227 1106 232
rect 1149 226 1152 232
rect 1203 226 1206 232
rect 1259 226 1262 232
rect 1313 226 1316 232
rect 1137 215 1140 223
rect 1137 211 1138 215
rect 1120 202 1123 205
rect 1137 189 1140 211
rect 1183 209 1186 222
rect 1183 206 1193 209
rect 1225 206 1228 210
rect 1237 212 1240 222
rect 1237 209 1256 212
rect 1285 212 1288 213
rect 1152 202 1154 205
rect 1174 202 1175 205
rect 1183 197 1186 206
rect 1150 194 1186 197
rect 1150 189 1153 194
rect 1183 189 1186 194
rect 1190 197 1193 206
rect 1204 202 1208 204
rect 1225 203 1229 206
rect 1204 201 1211 202
rect 1237 197 1240 209
rect 1287 208 1288 212
rect 1285 206 1288 208
rect 1261 202 1264 205
rect 1293 202 1296 222
rect 1319 215 1320 219
rect 1317 206 1320 215
rect 1347 211 1350 222
rect 1317 203 1318 206
rect 1336 202 1339 204
rect 1336 201 1342 202
rect 1293 197 1296 198
rect 1347 197 1350 207
rect 1204 194 1240 197
rect 1204 189 1207 194
rect 1237 189 1240 194
rect 1260 194 1296 197
rect 1260 189 1263 194
rect 1293 189 1296 194
rect 1314 194 1350 197
rect 1314 189 1317 194
rect 1347 189 1350 194
rect 1103 168 1106 185
rect 1166 168 1169 185
rect 1176 168 1179 171
rect 1220 168 1223 185
rect 1230 168 1233 171
rect 1276 168 1279 185
rect 1286 168 1289 171
rect 1330 168 1333 185
rect 1340 168 1343 171
rect 1361 168 1366 307
rect 999 165 1366 168
rect 1015 146 1018 165
rect 1098 163 1366 165
rect 1049 158 1050 161
rect 1049 131 1052 158
rect 1060 148 1064 150
rect 1098 146 1101 163
rect 1109 154 1141 157
rect 1043 127 1046 130
rect 1050 128 1052 131
rect 1060 131 1064 142
rect 1060 121 1063 131
rect 1115 126 1118 129
rect 1060 117 1061 121
rect 1132 120 1135 142
rect 1138 130 1141 154
rect 1161 146 1164 163
rect 1171 160 1174 163
rect 1215 146 1218 163
rect 1225 160 1228 163
rect 1271 146 1274 163
rect 1281 160 1284 163
rect 1325 146 1328 163
rect 1335 160 1338 163
rect 1145 137 1148 142
rect 1178 137 1181 142
rect 1145 134 1181 137
rect 1138 127 1143 130
rect 1147 126 1149 129
rect 1169 126 1170 129
rect 1178 125 1181 134
rect 1199 137 1202 142
rect 1232 137 1235 142
rect 1199 134 1235 137
rect 1255 137 1258 142
rect 1288 137 1291 142
rect 1255 134 1291 137
rect 1309 137 1312 142
rect 1342 137 1345 142
rect 1309 134 1345 137
rect 1185 125 1188 134
rect 1199 129 1206 130
rect 1199 127 1203 129
rect 1220 125 1224 128
rect 1178 122 1188 125
rect 1060 109 1063 117
rect 1132 116 1133 120
rect 1132 108 1135 116
rect 1178 109 1181 122
rect 1220 121 1223 125
rect 1232 122 1235 134
rect 1288 133 1291 134
rect 1256 126 1259 129
rect 1232 119 1251 122
rect 1232 109 1235 119
rect 1280 123 1283 125
rect 1268 115 1271 121
rect 1282 119 1283 123
rect 1280 118 1283 119
rect 1245 112 1271 115
rect 1288 109 1291 129
rect 1312 125 1313 128
rect 1331 129 1337 130
rect 1331 127 1334 129
rect 1312 116 1315 125
rect 1342 124 1345 134
rect 1314 112 1315 116
rect 1342 109 1345 120
rect 1026 99 1029 105
rect 1098 99 1101 104
rect 1144 99 1147 105
rect 1198 99 1201 105
rect 1254 99 1257 105
rect 1308 99 1311 105
rect 802 95 803 98
rect 780 94 803 95
rect 807 95 808 98
rect 986 96 1347 99
rect 807 94 814 95
rect 780 91 814 94
rect 818 91 824 95
rect 1170 93 1175 96
rect 1276 93 1280 96
rect 780 90 824 91
rect 656 87 824 90
rect 1102 90 1351 93
rect 656 86 780 87
rect 329 83 453 84
rect 442 76 446 83
rect 325 74 369 76
rect 418 74 462 76
rect 505 74 549 76
rect 325 72 549 74
rect 325 68 331 72
rect 335 71 424 72
rect 335 68 369 71
rect 418 68 424 71
rect 428 71 511 72
rect 428 68 462 71
rect 505 68 511 71
rect 515 68 549 72
rect 339 60 345 68
rect 339 56 340 60
rect 344 56 345 60
rect 350 62 354 63
rect 359 62 365 68
rect 400 62 411 65
rect 359 58 360 62
rect 364 58 365 62
rect 329 55 334 56
rect 329 51 330 55
rect 350 55 354 58
rect 329 48 334 51
rect 329 44 330 48
rect 329 43 334 44
rect 337 51 350 53
rect 337 49 354 51
rect 361 51 392 55
rect 329 42 333 43
rect 293 38 333 42
rect 329 25 333 38
rect 337 38 341 49
rect 352 42 357 46
rect 361 42 365 51
rect 344 34 347 38
rect 351 34 358 38
rect 337 30 341 34
rect 337 26 349 30
rect 353 29 358 34
rect 329 24 334 25
rect 329 20 330 24
rect 334 20 341 23
rect 329 17 341 20
rect 345 22 349 26
rect 352 25 368 29
rect 345 18 360 22
rect 364 18 365 22
rect 388 18 392 51
rect 408 52 411 62
rect 432 60 438 68
rect 432 56 433 60
rect 437 56 438 60
rect 443 62 447 63
rect 452 62 458 68
rect 452 58 453 62
rect 457 58 458 62
rect 519 60 525 68
rect 498 59 514 60
rect 422 55 427 56
rect 422 52 423 55
rect 408 51 423 52
rect 443 55 447 58
rect 408 49 427 51
rect 422 48 427 49
rect 422 44 423 48
rect 422 43 427 44
rect 430 51 443 53
rect 430 49 447 51
rect 422 25 426 43
rect 430 38 434 49
rect 454 46 458 55
rect 502 55 514 59
rect 519 56 520 60
rect 524 56 525 60
rect 530 62 534 63
rect 539 62 545 68
rect 539 58 540 62
rect 544 58 545 62
rect 502 54 510 55
rect 509 51 510 54
rect 530 55 534 58
rect 509 48 514 51
rect 445 42 450 46
rect 454 42 465 46
rect 509 44 510 48
rect 509 43 514 44
rect 517 51 530 53
rect 517 49 534 51
rect 437 34 440 38
rect 444 34 451 38
rect 430 30 434 34
rect 430 26 442 30
rect 422 24 427 25
rect 422 20 423 24
rect 427 20 434 23
rect 422 17 434 20
rect 438 22 442 26
rect 446 29 451 34
rect 446 25 461 29
rect 509 25 513 43
rect 517 38 521 49
rect 541 46 545 55
rect 532 42 537 46
rect 541 42 554 46
rect 524 34 527 38
rect 531 34 538 38
rect 517 30 521 34
rect 517 26 529 30
rect 509 24 514 25
rect 438 18 453 22
rect 457 18 458 22
rect 509 20 510 24
rect 514 20 521 23
rect 509 17 521 20
rect 525 22 529 26
rect 533 28 538 34
rect 533 25 546 28
rect 1000 29 1003 84
rect 1102 85 1105 90
rect 1148 84 1151 90
rect 1202 84 1205 90
rect 1258 84 1261 90
rect 1312 84 1315 90
rect 1136 73 1139 81
rect 1136 69 1137 73
rect 1119 60 1122 63
rect 1136 47 1139 69
rect 1182 67 1185 80
rect 1182 64 1192 67
rect 1224 64 1227 68
rect 1236 70 1239 80
rect 1236 67 1255 70
rect 1284 70 1287 71
rect 1151 60 1153 63
rect 1173 60 1174 63
rect 1182 55 1185 64
rect 1149 52 1185 55
rect 1149 47 1152 52
rect 1182 47 1185 52
rect 1189 55 1192 64
rect 1203 60 1207 62
rect 1224 61 1228 64
rect 1203 59 1210 60
rect 1236 55 1239 67
rect 1286 66 1287 70
rect 1284 64 1287 66
rect 1260 60 1263 63
rect 1292 60 1295 80
rect 1318 73 1319 77
rect 1316 64 1319 73
rect 1346 69 1349 80
rect 1316 61 1317 64
rect 1335 60 1338 62
rect 1335 59 1341 60
rect 1292 55 1295 56
rect 1346 55 1349 65
rect 1203 52 1239 55
rect 1203 47 1206 52
rect 1236 47 1239 52
rect 1259 52 1295 55
rect 1259 47 1262 52
rect 1292 47 1295 52
rect 1313 52 1349 55
rect 1313 47 1316 52
rect 1346 47 1349 52
rect 551 25 1005 29
rect 1000 24 1003 25
rect 1102 24 1105 43
rect 1165 24 1168 43
rect 1175 24 1178 29
rect 1219 24 1222 43
rect 1229 24 1232 29
rect 1275 24 1278 43
rect 1285 24 1288 29
rect 1329 24 1332 43
rect 1339 24 1342 29
rect 1360 24 1365 163
rect 525 18 540 22
rect 544 18 545 22
rect 1100 21 1365 24
rect 325 8 331 12
rect 335 8 341 12
rect 345 8 369 12
rect 418 8 424 12
rect 428 8 434 12
rect 438 8 462 12
rect 319 7 462 8
rect 505 8 511 12
rect 515 8 521 12
rect 525 8 549 12
rect 505 7 549 8
rect 319 5 549 7
rect 325 4 369 5
rect 418 4 549 5
<< metal2 >>
rect 363 455 468 456
rect 363 453 463 455
rect 81 448 110 452
rect 17 444 84 448
rect 17 302 22 444
rect 91 437 344 441
rect 32 379 36 430
rect 91 402 96 437
rect 339 433 343 437
rect 109 424 110 427
rect 114 424 198 427
rect 202 424 291 427
rect 295 424 316 427
rect 313 421 316 424
rect 363 421 367 453
rect 467 453 468 455
rect 474 423 478 457
rect 945 450 946 455
rect 516 438 764 442
rect 516 434 520 438
rect 573 426 662 429
rect 571 425 662 426
rect 666 425 749 429
rect 313 417 367 421
rect 195 406 339 409
rect 521 408 668 411
rect 90 398 102 402
rect 195 402 198 406
rect 665 404 668 408
rect 107 398 118 402
rect 247 397 248 400
rect 31 377 36 379
rect 31 341 35 377
rect 175 376 223 379
rect 175 375 232 376
rect 220 372 232 375
rect 245 366 248 397
rect 288 392 291 398
rect 569 400 573 403
rect 288 389 339 392
rect 569 392 572 400
rect 521 389 572 392
rect 665 400 666 404
rect 683 402 702 406
rect 760 404 764 438
rect 945 414 949 450
rect 1003 441 1025 444
rect 981 414 984 437
rect 1090 424 1170 427
rect 1090 418 1093 424
rect 1051 415 1093 418
rect 1166 418 1169 424
rect 1190 422 1249 425
rect 981 411 996 414
rect 1123 414 1144 417
rect 746 400 754 404
rect 759 402 764 404
rect 759 400 986 402
rect 566 381 569 389
rect 493 378 504 380
rect 566 378 580 381
rect 493 377 498 378
rect 274 374 498 377
rect 502 374 504 378
rect 274 373 504 374
rect 604 372 607 399
rect 666 390 669 400
rect 760 399 986 400
rect 773 398 986 399
rect 972 390 976 391
rect 666 386 976 390
rect 619 378 678 381
rect 509 369 607 372
rect 706 378 968 381
rect 692 374 696 377
rect 692 371 759 374
rect 197 365 250 366
rect 115 362 250 365
rect 509 364 513 369
rect 115 356 118 362
rect 64 353 129 356
rect 31 337 72 341
rect 68 330 72 337
rect 21 298 22 302
rect 29 328 32 329
rect 29 325 36 328
rect 29 260 32 325
rect 72 326 105 329
rect 125 329 128 353
rect 207 353 292 356
rect 296 353 317 356
rect 393 355 458 358
rect 176 325 209 328
rect 189 321 192 325
rect 301 321 304 327
rect 189 318 304 321
rect 265 309 266 312
rect 263 261 266 309
rect 314 303 317 353
rect 454 352 458 355
rect 509 352 512 364
rect 755 361 759 371
rect 516 358 536 360
rect 516 357 532 358
rect 516 353 517 357
rect 521 354 532 357
rect 536 355 621 358
rect 720 358 785 361
rect 521 353 536 354
rect 516 352 524 353
rect 454 349 512 352
rect 358 327 365 330
rect 308 299 342 303
rect 302 298 342 299
rect 29 257 123 260
rect 133 258 276 261
rect 120 253 123 257
rect 271 227 302 231
rect 252 226 276 227
rect 209 223 276 226
rect 209 222 212 223
rect 153 219 212 222
rect 153 210 157 219
rect 63 207 157 210
rect 28 179 35 182
rect 28 114 31 179
rect 71 180 104 183
rect 124 183 127 207
rect 206 207 291 210
rect 85 145 88 180
rect 175 179 208 182
rect 188 175 191 179
rect 300 175 303 181
rect 188 172 303 175
rect 264 163 265 166
rect 185 147 188 163
rect 85 141 178 145
rect 184 144 251 147
rect 173 128 178 141
rect 173 124 246 128
rect 262 115 265 163
rect 315 159 318 298
rect 326 275 347 279
rect 358 262 361 327
rect 401 328 434 331
rect 454 331 457 349
rect 593 347 751 350
rect 419 279 423 328
rect 505 327 538 330
rect 518 323 521 327
rect 630 323 633 329
rect 518 320 633 323
rect 685 330 692 333
rect 594 311 595 314
rect 592 263 595 311
rect 635 301 669 305
rect 629 300 669 301
rect 645 272 673 275
rect 685 265 688 330
rect 728 331 761 334
rect 781 334 784 358
rect 863 358 948 361
rect 840 350 914 352
rect 840 349 918 350
rect 744 276 748 331
rect 832 330 865 333
rect 845 326 848 330
rect 957 326 960 332
rect 845 323 960 326
rect 753 289 756 314
rect 921 314 922 317
rect 770 277 829 280
rect 837 276 841 314
rect 919 266 922 314
rect 358 259 452 262
rect 462 260 605 263
rect 685 262 779 265
rect 789 263 932 266
rect 449 255 452 259
rect 776 258 779 262
rect 747 251 767 254
rect 747 249 750 251
rect 507 246 750 249
rect 764 250 767 251
rect 827 251 875 254
rect 764 246 766 250
rect 770 246 771 249
rect 507 230 510 246
rect 827 242 830 251
rect 758 240 830 242
rect 754 239 830 240
rect 836 233 841 236
rect 327 227 510 230
rect 536 229 841 233
rect 536 228 659 229
rect 537 212 542 228
rect 869 215 872 251
rect 392 209 457 212
rect 424 193 427 209
rect 357 181 364 184
rect 310 158 340 159
rect 310 153 339 158
rect 280 124 300 128
rect 28 111 122 114
rect 132 112 275 115
rect 119 107 122 111
rect 311 10 317 153
rect 338 128 342 129
rect 326 124 342 128
rect 338 103 342 124
rect 357 116 360 181
rect 400 182 433 185
rect 453 185 456 209
rect 535 209 620 212
rect 719 212 784 215
rect 415 135 418 182
rect 504 181 537 184
rect 517 177 520 181
rect 629 177 632 183
rect 517 174 632 177
rect 684 184 691 187
rect 424 169 427 170
rect 593 165 594 168
rect 424 143 427 165
rect 415 131 514 135
rect 591 117 594 165
rect 633 155 669 158
rect 607 131 666 136
rect 684 119 687 184
rect 727 185 760 188
rect 780 188 783 212
rect 862 212 947 215
rect 747 149 751 185
rect 831 184 864 187
rect 844 180 847 184
rect 956 180 959 186
rect 844 177 959 180
rect 920 168 921 171
rect 731 145 751 149
rect 747 144 751 145
rect 705 133 832 136
rect 838 133 839 136
rect 705 132 839 133
rect 918 120 921 168
rect 357 113 451 116
rect 461 114 604 117
rect 684 116 778 119
rect 788 117 931 120
rect 448 109 451 113
rect 775 112 778 116
rect 727 108 731 109
rect 338 99 415 103
rect 412 95 415 99
rect 495 98 497 103
rect 495 95 500 98
rect 396 66 400 91
rect 412 91 500 95
rect 412 90 415 91
rect 727 59 731 104
rect 965 98 968 378
rect 502 56 731 59
rect 502 55 727 56
rect 964 46 968 98
rect 469 42 503 46
rect 558 43 968 46
rect 964 42 968 43
rect 499 38 503 42
rect 499 35 568 38
rect 565 31 568 35
rect 972 31 976 386
rect 373 25 461 29
rect 466 25 546 28
rect 565 27 976 31
rect 983 17 986 398
rect 993 302 996 411
rect 1127 408 1130 414
rect 1170 414 1196 417
rect 1200 414 1201 417
rect 1246 416 1249 422
rect 1270 417 1289 420
rect 1246 413 1253 416
rect 1270 412 1273 417
rect 1293 418 1332 419
rect 1293 416 1328 418
rect 1120 407 1130 408
rect 1156 407 1175 410
rect 1066 404 1078 407
rect 1120 405 1122 407
rect 1075 340 1078 404
rect 1126 405 1130 407
rect 1138 404 1159 407
rect 1172 404 1220 407
rect 1283 407 1342 410
rect 1253 402 1256 405
rect 1163 387 1166 399
rect 1088 384 1166 387
rect 1253 399 1311 402
rect 1088 355 1091 384
rect 1242 380 1246 398
rect 1123 376 1246 380
rect 1123 350 1127 376
rect 1242 375 1246 376
rect 1257 361 1315 364
rect 1142 356 1224 359
rect 1257 358 1260 361
rect 1287 353 1346 356
rect 1127 346 1148 349
rect 1174 346 1200 349
rect 1204 346 1205 349
rect 1250 347 1257 350
rect 1170 340 1173 346
rect 1075 337 1173 340
rect 1250 341 1253 347
rect 1297 345 1332 347
rect 1297 344 1336 345
rect 1194 338 1253 341
rect 1089 317 1161 319
rect 1085 315 1161 317
rect 993 299 1108 302
rect 993 298 1006 299
rect 1157 282 1161 315
rect 1303 308 1306 344
rect 1303 305 1401 308
rect 1090 279 1170 282
rect 1090 273 1093 279
rect 1051 270 1093 273
rect 1166 272 1169 279
rect 1190 277 1249 280
rect 1051 228 1054 270
rect 1123 269 1144 272
rect 1170 269 1196 272
rect 1200 269 1201 272
rect 1246 271 1249 277
rect 1270 272 1289 275
rect 1246 268 1253 271
rect 1270 267 1273 272
rect 1293 273 1332 274
rect 1293 271 1328 273
rect 1066 259 1078 262
rect 1050 162 1054 228
rect 1075 195 1078 259
rect 1138 259 1220 262
rect 1283 262 1342 265
rect 1253 257 1256 260
rect 1253 254 1311 257
rect 1242 235 1246 253
rect 1123 231 1246 235
rect 1123 205 1127 231
rect 1242 230 1246 231
rect 1257 216 1315 219
rect 1142 211 1224 214
rect 1257 213 1260 216
rect 1287 208 1346 211
rect 1127 201 1148 204
rect 1174 201 1200 204
rect 1204 201 1205 204
rect 1250 202 1257 205
rect 1170 195 1173 201
rect 1075 192 1173 195
rect 1250 196 1253 202
rect 1297 200 1332 202
rect 1297 199 1336 200
rect 1194 193 1253 196
rect 1302 174 1305 199
rect 1302 171 1373 174
rect 999 154 1046 157
rect 1000 88 1003 154
rect 1043 153 1046 154
rect 1062 154 1105 157
rect 1109 154 1110 157
rect 1062 153 1065 154
rect 1043 150 1065 153
rect 1089 137 1169 140
rect 1089 131 1092 137
rect 1050 128 1092 131
rect 1165 130 1168 137
rect 1189 135 1248 138
rect 1122 127 1143 130
rect 1169 127 1195 130
rect 1199 127 1200 130
rect 1245 129 1248 135
rect 1269 130 1288 133
rect 1245 126 1252 129
rect 1269 125 1272 130
rect 1292 131 1331 132
rect 1292 129 1327 131
rect 1065 117 1077 120
rect 1074 53 1077 117
rect 1137 117 1219 120
rect 1282 120 1341 123
rect 1252 115 1255 118
rect 1252 112 1310 115
rect 1241 93 1245 111
rect 1122 89 1245 93
rect 1122 63 1126 89
rect 1241 88 1245 89
rect 1256 74 1314 77
rect 1141 69 1223 72
rect 1256 71 1259 74
rect 1286 66 1345 69
rect 1126 59 1147 62
rect 1173 59 1199 62
rect 1203 59 1204 62
rect 1249 60 1256 63
rect 1169 53 1172 59
rect 1074 50 1172 53
rect 1249 54 1252 60
rect 1296 58 1331 60
rect 1296 57 1335 58
rect 1193 51 1252 54
rect 1302 29 1305 57
rect 1302 26 1370 29
rect 392 14 986 17
rect 311 3 312 10
<< metal3 >>
rect 497 378 522 380
rect 497 374 498 378
rect 502 374 522 378
rect 497 373 503 374
rect 516 359 522 374
rect 516 357 523 359
rect 516 353 517 357
rect 521 353 523 357
rect 516 352 523 353
<< ntransistor >>
rect 121 425 123 436
rect 128 425 130 436
rect 141 425 143 434
rect 208 425 210 436
rect 215 425 217 436
rect 228 425 230 434
rect 301 425 303 436
rect 308 425 310 436
rect 321 425 323 434
rect 541 427 543 436
rect 554 427 556 438
rect 561 427 563 438
rect 634 427 636 436
rect 647 427 649 438
rect 654 427 656 438
rect 721 427 723 436
rect 734 427 736 438
rect 741 427 743 438
rect 1042 392 1044 395
rect 1114 391 1116 394
rect 1153 391 1155 397
rect 1174 391 1176 397
rect 1207 391 1209 397
rect 1228 391 1230 397
rect 1263 391 1265 397
rect 1284 391 1286 397
rect 1317 391 1319 397
rect 1338 391 1340 397
rect 43 313 45 319
rect 55 307 57 316
rect 62 307 64 316
rect 121 315 123 324
rect 137 310 139 319
rect 147 310 149 319
rect 157 307 159 319
rect 164 307 166 319
rect 205 315 207 324
rect 221 310 223 319
rect 231 310 233 319
rect 241 307 243 319
rect 248 307 250 319
rect 275 313 277 319
rect 287 307 289 316
rect 294 307 296 316
rect 372 315 374 321
rect 384 309 386 318
rect 391 309 393 318
rect 450 317 452 326
rect 466 312 468 321
rect 476 312 478 321
rect 486 309 488 321
rect 493 309 495 321
rect 534 317 536 326
rect 550 312 552 321
rect 560 312 562 321
rect 570 309 572 321
rect 577 309 579 321
rect 604 315 606 321
rect 699 318 701 324
rect 1118 369 1120 372
rect 1157 366 1159 372
rect 1178 366 1180 372
rect 1211 366 1213 372
rect 1232 366 1234 372
rect 1267 366 1269 372
rect 1288 366 1290 372
rect 1321 366 1323 372
rect 1342 366 1344 372
rect 616 309 618 318
rect 623 309 625 318
rect 711 312 713 321
rect 718 312 720 321
rect 777 320 779 329
rect 793 315 795 324
rect 803 315 805 324
rect 813 312 815 324
rect 820 312 822 324
rect 861 320 863 329
rect 877 315 879 324
rect 887 315 889 324
rect 897 312 899 324
rect 904 312 906 324
rect 931 318 933 324
rect 943 312 945 321
rect 950 312 952 321
rect 136 279 138 285
rect 146 279 148 285
rect 156 279 158 285
rect 465 281 467 287
rect 475 281 477 287
rect 485 281 487 287
rect 792 284 794 290
rect 802 284 804 290
rect 812 284 814 290
rect 1042 247 1044 250
rect 1114 246 1116 249
rect 1153 246 1155 252
rect 1174 246 1176 252
rect 1207 246 1209 252
rect 1228 246 1230 252
rect 1263 246 1265 252
rect 1284 246 1286 252
rect 1317 246 1319 252
rect 1338 246 1340 252
rect 42 167 44 173
rect 54 161 56 170
rect 61 161 63 170
rect 120 169 122 178
rect 136 164 138 173
rect 146 164 148 173
rect 156 161 158 173
rect 163 161 165 173
rect 204 169 206 178
rect 220 164 222 173
rect 230 164 232 173
rect 240 161 242 173
rect 247 161 249 173
rect 274 167 276 173
rect 286 161 288 170
rect 293 161 295 170
rect 371 169 373 175
rect 383 163 385 172
rect 390 163 392 172
rect 449 171 451 180
rect 465 166 467 175
rect 475 166 477 175
rect 485 163 487 175
rect 492 163 494 175
rect 533 171 535 180
rect 549 166 551 175
rect 559 166 561 175
rect 569 163 571 175
rect 576 163 578 175
rect 603 169 605 175
rect 698 172 700 178
rect 1118 224 1120 227
rect 1157 221 1159 227
rect 1178 221 1180 227
rect 1211 221 1213 227
rect 1232 221 1234 227
rect 1267 221 1269 227
rect 1288 221 1290 227
rect 1321 221 1323 227
rect 1342 221 1344 227
rect 615 163 617 172
rect 622 163 624 172
rect 710 166 712 175
rect 717 166 719 175
rect 776 174 778 183
rect 792 169 794 178
rect 802 169 804 178
rect 812 166 814 178
rect 819 166 821 178
rect 860 174 862 183
rect 876 169 878 178
rect 886 169 888 178
rect 896 166 898 178
rect 903 166 905 178
rect 930 172 932 178
rect 942 166 944 175
rect 949 166 951 175
rect 135 133 137 139
rect 145 133 147 139
rect 155 133 157 139
rect 464 135 466 141
rect 474 135 476 141
rect 484 135 486 141
rect 791 138 793 144
rect 801 138 803 144
rect 811 138 813 144
rect 1041 105 1043 108
rect 1113 104 1115 107
rect 1152 104 1154 110
rect 1173 104 1175 110
rect 1206 104 1208 110
rect 1227 104 1229 110
rect 1262 104 1264 110
rect 1283 104 1285 110
rect 1316 104 1318 110
rect 1337 104 1339 110
rect 1117 82 1119 85
rect 1156 79 1158 85
rect 1177 79 1179 85
rect 1210 79 1212 85
rect 1231 79 1233 85
rect 1266 79 1268 85
rect 1287 79 1289 85
rect 1320 79 1322 85
rect 1341 79 1343 85
rect 336 19 338 28
rect 349 17 351 28
rect 356 17 358 28
rect 429 19 431 28
rect 442 17 444 28
rect 449 17 451 28
rect 516 19 518 28
rect 529 17 531 28
rect 536 17 538 28
<< ptransistor >>
rect 1042 428 1044 434
rect 1114 428 1116 434
rect 1153 428 1155 434
rect 1174 428 1176 434
rect 1207 428 1209 434
rect 1228 428 1230 434
rect 1263 428 1265 434
rect 1284 428 1286 434
rect 1317 428 1319 434
rect 1338 428 1340 434
rect 121 390 123 403
rect 131 390 133 403
rect 141 392 143 410
rect 208 390 210 403
rect 218 390 220 403
rect 228 392 230 410
rect 301 390 303 403
rect 311 390 313 403
rect 321 392 323 410
rect 541 394 543 412
rect 551 392 553 405
rect 561 392 563 405
rect 634 394 636 412
rect 644 392 646 405
rect 654 392 656 405
rect 721 394 723 412
rect 731 392 733 405
rect 741 392 743 405
rect 43 336 45 348
rect 53 336 55 346
rect 63 336 65 346
rect 129 337 131 364
rect 145 337 147 355
rect 155 337 157 355
rect 165 337 167 364
rect 213 337 215 364
rect 229 337 231 355
rect 239 337 241 355
rect 249 337 251 364
rect 275 336 277 348
rect 285 336 287 346
rect 295 336 297 346
rect 372 338 374 350
rect 382 338 384 348
rect 392 338 394 348
rect 458 339 460 366
rect 474 339 476 357
rect 484 339 486 357
rect 494 339 496 366
rect 542 339 544 366
rect 558 339 560 357
rect 568 339 570 357
rect 578 339 580 366
rect 604 338 606 350
rect 614 338 616 348
rect 624 338 626 348
rect 699 341 701 353
rect 709 341 711 351
rect 719 341 721 351
rect 785 342 787 369
rect 801 342 803 360
rect 811 342 813 360
rect 821 342 823 369
rect 869 342 871 369
rect 885 342 887 360
rect 895 342 897 360
rect 905 342 907 369
rect 931 341 933 353
rect 941 341 943 351
rect 951 341 953 351
rect 1118 329 1120 335
rect 1157 329 1159 335
rect 1178 329 1180 335
rect 1211 329 1213 335
rect 1232 329 1234 335
rect 1267 329 1269 335
rect 1288 329 1290 335
rect 1321 329 1323 335
rect 1342 329 1344 335
rect 136 234 138 252
rect 143 234 145 252
rect 156 243 158 255
rect 1042 283 1044 289
rect 1114 283 1116 289
rect 1153 283 1155 289
rect 1174 283 1176 289
rect 1207 283 1209 289
rect 1228 283 1230 289
rect 1263 283 1265 289
rect 1284 283 1286 289
rect 1317 283 1319 289
rect 1338 283 1340 289
rect 465 236 467 254
rect 472 236 474 254
rect 485 245 487 257
rect 792 239 794 257
rect 799 239 801 257
rect 812 248 814 260
rect 42 190 44 202
rect 52 190 54 200
rect 62 190 64 200
rect 128 191 130 218
rect 144 191 146 209
rect 154 191 156 209
rect 164 191 166 218
rect 212 191 214 218
rect 228 191 230 209
rect 238 191 240 209
rect 248 191 250 218
rect 274 190 276 202
rect 284 190 286 200
rect 294 190 296 200
rect 371 192 373 204
rect 381 192 383 202
rect 391 192 393 202
rect 457 193 459 220
rect 473 193 475 211
rect 483 193 485 211
rect 493 193 495 220
rect 541 193 543 220
rect 557 193 559 211
rect 567 193 569 211
rect 577 193 579 220
rect 603 192 605 204
rect 613 192 615 202
rect 623 192 625 202
rect 698 195 700 207
rect 708 195 710 205
rect 718 195 720 205
rect 784 196 786 223
rect 800 196 802 214
rect 810 196 812 214
rect 820 196 822 223
rect 868 196 870 223
rect 884 196 886 214
rect 894 196 896 214
rect 904 196 906 223
rect 930 195 932 207
rect 940 195 942 205
rect 950 195 952 205
rect 1118 184 1120 190
rect 1157 184 1159 190
rect 1178 184 1180 190
rect 1211 184 1213 190
rect 1232 184 1234 190
rect 1267 184 1269 190
rect 1288 184 1290 190
rect 1321 184 1323 190
rect 1342 184 1344 190
rect 1041 141 1043 147
rect 1113 141 1115 147
rect 1152 141 1154 147
rect 1173 141 1175 147
rect 1206 141 1208 147
rect 1227 141 1229 147
rect 1262 141 1264 147
rect 1283 141 1285 147
rect 1316 141 1318 147
rect 1337 141 1339 147
rect 135 88 137 106
rect 142 88 144 106
rect 155 97 157 109
rect 464 90 466 108
rect 471 90 473 108
rect 484 99 486 111
rect 791 93 793 111
rect 798 93 800 111
rect 811 102 813 114
rect 336 43 338 61
rect 346 50 348 63
rect 356 50 358 63
rect 429 43 431 61
rect 439 50 441 63
rect 449 50 451 63
rect 516 43 518 61
rect 526 50 528 63
rect 536 50 538 63
rect 1117 42 1119 48
rect 1156 42 1158 48
rect 1177 42 1179 48
rect 1210 42 1212 48
rect 1231 42 1233 48
rect 1266 42 1268 48
rect 1287 42 1289 48
rect 1320 42 1322 48
rect 1341 42 1343 48
<< polycontact >>
rect 128 415 132 419
rect 138 415 142 419
rect 118 407 122 411
rect 215 415 219 419
rect 225 415 229 419
rect 205 407 209 411
rect 308 415 312 419
rect 318 415 322 419
rect 298 407 302 411
rect 542 417 546 421
rect 552 417 556 421
rect 635 417 639 421
rect 645 417 649 421
rect 562 409 566 413
rect 722 417 726 421
rect 732 417 736 421
rect 655 409 659 413
rect 1040 413 1044 417
rect 742 409 746 413
rect 1112 412 1116 416
rect 1150 412 1154 416
rect 1171 412 1175 416
rect 1204 412 1208 416
rect 1225 412 1229 416
rect 1260 412 1264 416
rect 1281 412 1285 416
rect 1314 412 1318 416
rect 1335 412 1339 416
rect 54 352 58 356
rect 115 344 119 348
rect 44 328 48 332
rect 199 344 203 348
rect 152 329 156 333
rect 162 329 166 333
rect 286 352 290 356
rect 383 354 387 358
rect 444 346 448 350
rect 63 320 67 324
rect 131 323 135 327
rect 236 329 240 333
rect 246 329 250 333
rect 276 328 280 332
rect 215 323 219 327
rect 373 330 377 334
rect 295 320 299 324
rect 528 346 532 350
rect 481 331 485 335
rect 491 331 495 335
rect 615 354 619 358
rect 710 357 714 361
rect 771 349 775 353
rect 392 322 396 326
rect 460 325 464 329
rect 565 331 569 335
rect 575 331 579 335
rect 605 330 609 334
rect 544 325 548 329
rect 700 333 704 337
rect 624 322 628 326
rect 855 349 859 353
rect 808 334 812 338
rect 818 334 822 338
rect 942 357 946 361
rect 1116 347 1120 351
rect 1154 347 1158 351
rect 1175 347 1179 351
rect 1208 347 1212 351
rect 1229 347 1233 351
rect 1264 347 1268 351
rect 1285 347 1289 351
rect 1318 347 1322 351
rect 1339 347 1343 351
rect 719 325 723 329
rect 787 328 791 332
rect 892 334 896 338
rect 902 334 906 338
rect 932 333 936 337
rect 871 328 875 332
rect 951 325 955 329
rect 133 266 137 270
rect 145 266 149 270
rect 153 265 157 269
rect 462 268 466 272
rect 474 268 478 272
rect 143 258 147 262
rect 482 267 486 271
rect 789 271 793 275
rect 801 271 805 275
rect 472 260 476 264
rect 809 270 813 274
rect 799 263 803 267
rect 1040 268 1044 272
rect 1112 267 1116 271
rect 1150 267 1154 271
rect 1171 267 1175 271
rect 1204 267 1208 271
rect 1225 267 1229 271
rect 1260 267 1264 271
rect 1281 267 1285 271
rect 1314 267 1318 271
rect 1335 267 1339 271
rect 53 206 57 210
rect 114 198 118 202
rect 43 182 47 186
rect 198 198 202 202
rect 151 183 155 187
rect 161 183 165 187
rect 285 206 289 210
rect 382 208 386 212
rect 443 200 447 204
rect 62 174 66 178
rect 130 177 134 181
rect 235 183 239 187
rect 245 183 249 187
rect 275 182 279 186
rect 214 177 218 181
rect 372 184 376 188
rect 294 174 298 178
rect 527 200 531 204
rect 480 185 484 189
rect 490 185 494 189
rect 614 208 618 212
rect 709 211 713 215
rect 770 203 774 207
rect 391 176 395 180
rect 459 179 463 183
rect 564 185 568 189
rect 574 185 578 189
rect 604 184 608 188
rect 543 179 547 183
rect 699 187 703 191
rect 623 176 627 180
rect 854 203 858 207
rect 807 188 811 192
rect 817 188 821 192
rect 941 211 945 215
rect 1116 202 1120 206
rect 1154 202 1158 206
rect 1175 202 1179 206
rect 1208 202 1212 206
rect 1229 202 1233 206
rect 1264 202 1268 206
rect 1285 202 1289 206
rect 1318 202 1322 206
rect 1339 202 1343 206
rect 718 179 722 183
rect 786 182 790 186
rect 891 188 895 192
rect 901 188 905 192
rect 931 187 935 191
rect 870 182 874 186
rect 950 179 954 183
rect 132 120 136 124
rect 144 120 148 124
rect 152 119 156 123
rect 461 122 465 126
rect 473 122 477 126
rect 142 112 146 116
rect 481 121 485 125
rect 788 125 792 129
rect 800 125 804 129
rect 471 114 475 118
rect 808 124 812 128
rect 1039 126 1043 130
rect 798 117 802 121
rect 1111 125 1115 129
rect 1149 125 1153 129
rect 1170 125 1174 129
rect 1203 125 1207 129
rect 1224 125 1228 129
rect 1259 125 1263 129
rect 1280 125 1284 129
rect 1313 125 1317 129
rect 1334 125 1338 129
rect 357 42 361 46
rect 337 34 341 38
rect 347 34 351 38
rect 450 42 454 46
rect 1115 60 1119 64
rect 1153 60 1157 64
rect 1174 60 1178 64
rect 1207 60 1211 64
rect 1228 60 1232 64
rect 1263 60 1267 64
rect 1284 60 1288 64
rect 1317 60 1321 64
rect 1338 60 1342 64
rect 430 34 434 38
rect 440 34 444 38
rect 537 42 541 46
rect 517 34 521 38
rect 527 34 531 38
<< ndcontact >>
rect 134 441 138 445
rect 221 441 225 445
rect 115 431 119 435
rect 314 441 318 445
rect 145 429 149 433
rect 202 431 206 435
rect 546 443 550 447
rect 232 429 236 433
rect 295 431 299 435
rect 639 443 643 447
rect 325 429 329 433
rect 535 431 539 435
rect 565 433 569 437
rect 726 443 730 447
rect 628 431 632 435
rect 658 433 662 437
rect 715 431 719 435
rect 745 433 749 437
rect 1027 392 1031 396
rect 1061 392 1065 396
rect 1099 391 1103 395
rect 1133 391 1137 395
rect 1145 392 1149 396
rect 1179 392 1183 396
rect 1199 392 1203 396
rect 1233 392 1237 396
rect 1255 392 1259 396
rect 1289 392 1293 396
rect 1309 392 1313 396
rect 1343 392 1347 396
rect 37 314 41 318
rect 115 319 119 323
rect 199 319 203 323
rect 66 311 70 315
rect 129 311 133 315
rect 141 314 145 318
rect 151 312 155 316
rect 48 302 52 306
rect 213 311 217 315
rect 225 314 229 318
rect 235 312 239 316
rect 169 302 173 306
rect 269 314 273 318
rect 366 316 370 320
rect 444 321 448 325
rect 298 311 302 315
rect 528 321 532 325
rect 395 313 399 317
rect 458 313 462 317
rect 470 316 474 320
rect 480 314 484 318
rect 253 302 257 306
rect 280 302 284 306
rect 377 304 381 308
rect 542 313 546 317
rect 554 316 558 320
rect 564 314 568 318
rect 498 304 502 308
rect 598 316 602 320
rect 693 319 697 323
rect 1103 368 1107 372
rect 1137 368 1141 372
rect 1149 367 1153 371
rect 1183 367 1187 371
rect 1203 367 1207 371
rect 1237 367 1241 371
rect 1259 367 1263 371
rect 1293 367 1297 371
rect 1313 367 1317 371
rect 1347 367 1351 371
rect 771 324 775 328
rect 627 313 631 317
rect 855 324 859 328
rect 722 316 726 320
rect 785 316 789 320
rect 797 319 801 323
rect 807 317 811 321
rect 582 304 586 308
rect 609 304 613 308
rect 704 307 708 311
rect 869 316 873 320
rect 881 319 885 323
rect 891 317 895 321
rect 825 307 829 311
rect 925 319 929 323
rect 954 316 958 320
rect 909 307 913 311
rect 936 307 940 311
rect 130 280 134 284
rect 140 280 144 284
rect 150 280 154 284
rect 160 280 164 284
rect 459 282 463 286
rect 469 282 473 286
rect 479 282 483 286
rect 489 282 493 286
rect 786 285 790 289
rect 796 285 800 289
rect 806 285 810 289
rect 816 285 820 289
rect 1027 247 1031 251
rect 1061 247 1065 251
rect 1099 246 1103 250
rect 1133 246 1137 250
rect 1145 247 1149 251
rect 1179 247 1183 251
rect 1199 247 1203 251
rect 1233 247 1237 251
rect 1255 247 1259 251
rect 1289 247 1293 251
rect 1309 247 1313 251
rect 1343 247 1347 251
rect 36 168 40 172
rect 114 173 118 177
rect 198 173 202 177
rect 65 165 69 169
rect 128 165 132 169
rect 140 168 144 172
rect 150 166 154 170
rect 47 156 51 160
rect 212 165 216 169
rect 224 168 228 172
rect 234 166 238 170
rect 168 156 172 160
rect 268 168 272 172
rect 365 170 369 174
rect 443 175 447 179
rect 297 165 301 169
rect 527 175 531 179
rect 394 167 398 171
rect 457 167 461 171
rect 469 170 473 174
rect 479 168 483 172
rect 252 156 256 160
rect 279 156 283 160
rect 376 158 380 162
rect 541 167 545 171
rect 553 170 557 174
rect 563 168 567 172
rect 497 158 501 162
rect 597 170 601 174
rect 692 173 696 177
rect 1103 223 1107 227
rect 1137 223 1141 227
rect 1149 222 1153 226
rect 1183 222 1187 226
rect 1203 222 1207 226
rect 1237 222 1241 226
rect 1259 222 1263 226
rect 1293 222 1297 226
rect 1313 222 1317 226
rect 1347 222 1351 226
rect 770 178 774 182
rect 626 167 630 171
rect 854 178 858 182
rect 721 170 725 174
rect 784 170 788 174
rect 796 173 800 177
rect 806 171 810 175
rect 581 158 585 162
rect 608 158 612 162
rect 703 161 707 165
rect 868 170 872 174
rect 880 173 884 177
rect 890 171 894 175
rect 824 161 828 165
rect 924 173 928 177
rect 953 170 957 174
rect 908 161 912 165
rect 935 161 939 165
rect 129 134 133 138
rect 139 134 143 138
rect 149 134 153 138
rect 159 134 163 138
rect 458 136 462 140
rect 468 136 472 140
rect 478 136 482 140
rect 488 136 492 140
rect 785 139 789 143
rect 795 139 799 143
rect 805 139 809 143
rect 815 139 819 143
rect 1026 105 1030 109
rect 1060 105 1064 109
rect 1098 104 1102 108
rect 1132 104 1136 108
rect 1144 105 1148 109
rect 1178 105 1182 109
rect 1198 105 1202 109
rect 1232 105 1236 109
rect 1254 105 1258 109
rect 1288 105 1292 109
rect 1308 105 1312 109
rect 1342 105 1346 109
rect 1102 81 1106 85
rect 1136 81 1140 85
rect 1148 80 1152 84
rect 1182 80 1186 84
rect 1202 80 1206 84
rect 1236 80 1240 84
rect 1258 80 1262 84
rect 1292 80 1296 84
rect 1312 80 1316 84
rect 1346 80 1350 84
rect 330 20 334 24
rect 360 18 364 22
rect 423 20 427 24
rect 453 18 457 22
rect 510 20 514 24
rect 341 8 345 12
rect 540 18 544 22
rect 434 8 438 12
rect 521 8 525 12
<< pdcontact >>
rect 1016 429 1020 433
rect 1060 429 1066 435
rect 1099 429 1103 433
rect 1132 429 1136 433
rect 1145 429 1149 433
rect 1162 429 1166 433
rect 1179 429 1183 433
rect 1199 429 1203 433
rect 1216 429 1220 433
rect 1233 429 1237 433
rect 1255 429 1259 433
rect 1272 429 1276 433
rect 1289 429 1293 433
rect 1309 429 1313 433
rect 1326 429 1330 433
rect 1343 429 1347 433
rect 115 391 119 395
rect 125 398 129 402
rect 125 391 129 395
rect 135 393 139 397
rect 145 405 149 409
rect 145 398 149 402
rect 202 391 206 395
rect 212 398 216 402
rect 212 391 216 395
rect 222 393 226 397
rect 232 405 236 409
rect 232 398 236 402
rect 295 391 299 395
rect 305 398 309 402
rect 305 391 309 395
rect 315 393 319 397
rect 325 405 329 409
rect 325 398 329 402
rect 535 407 539 411
rect 535 400 539 404
rect 628 407 632 411
rect 545 395 549 399
rect 555 400 559 404
rect 555 393 559 397
rect 628 400 632 404
rect 565 393 569 397
rect 715 407 719 411
rect 638 395 642 399
rect 648 400 652 404
rect 648 393 652 397
rect 715 400 719 404
rect 658 393 662 397
rect 725 395 729 399
rect 735 400 739 404
rect 735 393 739 397
rect 745 393 749 397
rect 37 337 41 341
rect 47 337 51 341
rect 57 337 61 341
rect 67 341 71 345
rect 123 338 127 342
rect 133 359 137 363
rect 133 352 137 356
rect 149 338 153 342
rect 159 345 163 349
rect 169 353 173 357
rect 207 338 211 342
rect 217 359 221 363
rect 217 352 221 356
rect 233 338 237 342
rect 243 345 247 349
rect 253 353 257 357
rect 269 337 273 341
rect 279 337 283 341
rect 289 337 293 341
rect 299 341 303 345
rect 366 339 370 343
rect 376 339 380 343
rect 386 339 390 343
rect 396 343 400 347
rect 452 340 456 344
rect 462 361 466 365
rect 462 354 466 358
rect 478 340 482 344
rect 488 347 492 351
rect 498 355 502 359
rect 536 340 540 344
rect 546 361 550 365
rect 546 354 550 358
rect 562 340 566 344
rect 572 347 576 351
rect 582 355 586 359
rect 598 339 602 343
rect 608 339 612 343
rect 618 339 622 343
rect 628 343 632 347
rect 693 342 697 346
rect 703 342 707 346
rect 713 342 717 346
rect 723 346 727 350
rect 779 343 783 347
rect 789 364 793 368
rect 789 357 793 361
rect 805 343 809 347
rect 815 350 819 354
rect 825 358 829 362
rect 863 343 867 347
rect 873 364 877 368
rect 873 357 877 361
rect 889 343 893 347
rect 899 350 903 354
rect 909 358 913 362
rect 925 342 929 346
rect 935 342 939 346
rect 945 342 949 346
rect 955 346 959 350
rect 1103 330 1107 334
rect 1136 330 1140 334
rect 1149 330 1153 334
rect 1166 330 1170 334
rect 1183 330 1187 334
rect 1203 330 1207 334
rect 1220 330 1224 334
rect 1237 330 1241 334
rect 1259 330 1263 334
rect 1276 330 1280 334
rect 1293 330 1297 334
rect 1313 330 1317 334
rect 1330 330 1334 334
rect 1347 330 1351 334
rect 1016 284 1020 288
rect 130 242 134 246
rect 1060 284 1066 290
rect 1099 284 1103 288
rect 1132 284 1136 288
rect 1145 284 1149 288
rect 1162 284 1166 288
rect 1179 284 1183 288
rect 1199 284 1203 288
rect 1216 284 1220 288
rect 1233 284 1237 288
rect 1255 284 1259 288
rect 1272 284 1276 288
rect 1289 284 1293 288
rect 1309 284 1313 288
rect 1326 284 1330 288
rect 1343 284 1347 288
rect 160 244 164 248
rect 459 244 463 248
rect 148 235 152 239
rect 489 246 493 250
rect 786 247 790 251
rect 477 237 481 241
rect 816 249 820 253
rect 804 240 808 244
rect 36 191 40 195
rect 46 191 50 195
rect 56 191 60 195
rect 66 195 70 199
rect 122 192 126 196
rect 132 213 136 217
rect 132 206 136 210
rect 148 192 152 196
rect 158 199 162 203
rect 168 207 172 211
rect 206 192 210 196
rect 216 213 220 217
rect 216 206 220 210
rect 232 192 236 196
rect 242 199 246 203
rect 252 207 256 211
rect 268 191 272 195
rect 278 191 282 195
rect 288 191 292 195
rect 298 195 302 199
rect 365 193 369 197
rect 375 193 379 197
rect 385 193 389 197
rect 395 197 399 201
rect 451 194 455 198
rect 461 215 465 219
rect 461 208 465 212
rect 477 194 481 198
rect 487 201 491 205
rect 497 209 501 213
rect 535 194 539 198
rect 545 215 549 219
rect 545 208 549 212
rect 561 194 565 198
rect 571 201 575 205
rect 581 209 585 213
rect 597 193 601 197
rect 607 193 611 197
rect 617 193 621 197
rect 627 197 631 201
rect 692 196 696 200
rect 702 196 706 200
rect 712 196 716 200
rect 722 200 726 204
rect 778 197 782 201
rect 788 218 792 222
rect 788 211 792 215
rect 804 197 808 201
rect 814 204 818 208
rect 824 212 828 216
rect 862 197 866 201
rect 872 218 876 222
rect 872 211 876 215
rect 888 197 892 201
rect 898 204 902 208
rect 908 212 912 216
rect 924 196 928 200
rect 934 196 938 200
rect 944 196 948 200
rect 954 200 958 204
rect 1103 185 1107 189
rect 1136 185 1140 189
rect 1149 185 1153 189
rect 1166 185 1170 189
rect 1183 185 1187 189
rect 1203 185 1207 189
rect 1220 185 1224 189
rect 1237 185 1241 189
rect 1259 185 1263 189
rect 1276 185 1280 189
rect 1293 185 1297 189
rect 1313 185 1317 189
rect 1330 185 1334 189
rect 1347 185 1351 189
rect 1015 142 1019 146
rect 1059 142 1065 148
rect 1098 142 1102 146
rect 1131 142 1135 146
rect 1144 142 1148 146
rect 1161 142 1165 146
rect 1178 142 1182 146
rect 1198 142 1202 146
rect 1215 142 1219 146
rect 1232 142 1236 146
rect 1254 142 1258 146
rect 1271 142 1275 146
rect 1288 142 1292 146
rect 1308 142 1312 146
rect 1325 142 1329 146
rect 1342 142 1346 146
rect 129 96 133 100
rect 159 98 163 102
rect 458 98 462 102
rect 147 89 151 93
rect 488 100 492 104
rect 785 101 789 105
rect 476 91 480 95
rect 815 103 819 107
rect 803 94 807 98
rect 330 51 334 55
rect 330 44 334 48
rect 340 56 344 60
rect 350 58 354 62
rect 350 51 354 55
rect 360 58 364 62
rect 423 51 427 55
rect 423 44 427 48
rect 433 56 437 60
rect 443 58 447 62
rect 443 51 447 55
rect 453 58 457 62
rect 510 51 514 55
rect 510 44 514 48
rect 520 56 524 60
rect 530 58 534 62
rect 530 51 534 55
rect 540 58 544 62
rect 1102 43 1106 47
rect 1135 43 1139 47
rect 1148 43 1152 47
rect 1165 43 1169 47
rect 1182 43 1186 47
rect 1202 43 1206 47
rect 1219 43 1223 47
rect 1236 43 1240 47
rect 1258 43 1262 47
rect 1275 43 1279 47
rect 1292 43 1296 47
rect 1312 43 1316 47
rect 1329 43 1333 47
rect 1346 43 1350 47
<< m2contact >>
rect 474 457 479 463
rect 110 448 115 453
rect 463 451 467 455
rect 946 450 951 455
rect 999 441 1003 445
rect 32 430 37 436
rect 110 424 114 428
rect 102 398 107 403
rect 198 424 202 428
rect 194 398 198 402
rect 291 424 295 428
rect 339 429 343 433
rect 515 429 520 434
rect 243 397 247 401
rect 287 398 291 402
rect 980 437 984 441
rect 473 418 478 423
rect 569 426 573 430
rect 339 406 343 410
rect 516 406 521 411
rect 573 400 577 404
rect 339 389 343 393
rect 517 389 521 393
rect 604 399 608 404
rect 662 425 666 429
rect 1025 441 1029 445
rect 749 425 753 429
rect 666 400 670 404
rect 679 402 683 406
rect 232 372 236 376
rect 269 373 274 377
rect 580 378 585 383
rect 615 378 619 383
rect 678 378 682 382
rect 692 377 696 381
rect 702 402 706 406
rect 944 408 950 414
rect 1047 414 1051 418
rect 1119 413 1123 417
rect 754 400 759 404
rect 702 378 706 382
rect 1062 404 1066 408
rect 1122 403 1126 407
rect 1144 413 1148 417
rect 1166 414 1170 418
rect 1134 403 1138 407
rect 1186 421 1190 425
rect 1196 413 1200 417
rect 1163 399 1167 403
rect 1220 404 1224 408
rect 1253 413 1257 417
rect 1289 416 1293 420
rect 1252 405 1256 409
rect 1269 408 1273 412
rect 1279 406 1283 410
rect 1242 398 1246 402
rect 1328 414 1332 418
rect 1342 407 1346 411
rect 1311 399 1315 403
rect 60 352 64 356
rect 203 352 207 356
rect 36 324 40 328
rect 68 326 72 330
rect 105 326 109 330
rect 125 325 129 329
rect 172 325 176 329
rect 209 325 213 329
rect 292 352 296 356
rect 261 309 265 313
rect 300 327 304 331
rect 17 298 21 302
rect 302 299 308 305
rect 129 257 133 261
rect 120 249 124 253
rect 322 275 326 279
rect 389 354 393 358
rect 532 354 536 358
rect 365 326 369 330
rect 397 328 401 332
rect 434 328 438 332
rect 454 327 458 331
rect 589 347 593 351
rect 501 327 505 331
rect 538 327 542 331
rect 621 354 625 358
rect 590 311 594 315
rect 629 329 633 333
rect 342 298 349 305
rect 629 301 635 307
rect 347 275 351 279
rect 419 275 423 279
rect 458 259 462 263
rect 449 251 453 255
rect 641 272 645 276
rect 716 357 720 361
rect 859 357 863 361
rect 751 347 755 351
rect 692 329 696 333
rect 724 331 728 335
rect 761 331 765 335
rect 781 330 785 334
rect 836 349 840 353
rect 828 330 832 334
rect 752 314 756 318
rect 837 314 841 318
rect 914 350 919 354
rect 865 330 869 334
rect 948 357 952 361
rect 917 314 921 318
rect 956 332 960 336
rect 1138 356 1142 360
rect 1086 350 1091 355
rect 669 300 676 307
rect 753 284 758 289
rect 673 272 677 276
rect 744 272 748 276
rect 302 227 307 231
rect 322 226 327 231
rect 766 277 770 281
rect 785 262 789 266
rect 776 254 780 258
rect 829 277 833 281
rect 837 271 841 276
rect 766 246 770 250
rect 754 240 758 244
rect 836 236 841 243
rect 1123 346 1127 350
rect 1224 355 1228 359
rect 1256 354 1260 358
rect 1148 346 1152 350
rect 1170 346 1174 350
rect 1200 346 1204 350
rect 1283 353 1287 357
rect 1257 346 1261 350
rect 1315 360 1319 364
rect 1346 352 1350 356
rect 1293 343 1297 347
rect 1332 345 1336 349
rect 1190 338 1194 342
rect 1084 317 1089 322
rect 1108 299 1112 303
rect 1047 269 1051 273
rect 1119 268 1123 272
rect 1062 259 1066 263
rect 1144 268 1148 272
rect 1166 268 1170 272
rect 1186 276 1190 280
rect 1196 268 1200 272
rect 1134 258 1138 262
rect 1220 259 1224 263
rect 1253 268 1257 272
rect 1289 271 1293 275
rect 1252 260 1256 264
rect 1269 263 1273 267
rect 1279 261 1283 265
rect 1242 253 1246 257
rect 1328 269 1332 273
rect 1342 262 1346 266
rect 1311 254 1315 258
rect 59 206 63 210
rect 35 178 39 182
rect 67 180 71 184
rect 104 180 108 184
rect 124 179 128 183
rect 171 179 175 183
rect 202 206 206 210
rect 208 179 212 183
rect 185 163 189 167
rect 291 206 295 210
rect 260 163 264 167
rect 299 181 303 185
rect 302 153 310 160
rect 251 143 255 147
rect 128 111 132 115
rect 119 103 123 107
rect 246 124 252 130
rect 275 124 280 129
rect 300 124 305 129
rect 321 124 326 129
rect 388 208 392 212
rect 531 208 535 212
rect 424 189 428 193
rect 364 180 368 184
rect 396 182 400 186
rect 433 182 437 186
rect 453 181 457 185
rect 500 181 504 185
rect 424 165 428 169
rect 537 181 541 185
rect 620 208 624 212
rect 589 165 593 169
rect 628 183 632 187
rect 339 153 344 158
rect 629 154 633 158
rect 424 139 428 143
rect 424 121 428 125
rect 457 113 461 117
rect 448 105 452 109
rect 514 131 520 136
rect 602 131 607 136
rect 715 211 719 215
rect 858 211 862 215
rect 691 183 695 187
rect 723 185 727 189
rect 760 185 764 189
rect 780 184 784 188
rect 827 184 831 188
rect 864 184 868 188
rect 947 211 951 215
rect 916 168 920 172
rect 955 186 959 190
rect 669 154 673 158
rect 727 145 731 149
rect 666 131 671 136
rect 700 131 705 136
rect 497 98 502 103
rect 396 91 400 95
rect 784 116 788 120
rect 775 108 779 112
rect 832 133 838 138
rect 727 104 731 108
rect 1138 211 1142 215
rect 1123 201 1127 205
rect 1224 210 1228 214
rect 1256 209 1260 213
rect 1148 201 1152 205
rect 1170 201 1174 205
rect 1200 201 1204 205
rect 1283 208 1287 212
rect 1257 201 1261 205
rect 1315 215 1319 219
rect 1346 207 1350 211
rect 1293 198 1297 202
rect 1332 200 1336 204
rect 1190 193 1194 197
rect 1050 158 1054 162
rect 1105 154 1109 158
rect 1046 127 1050 131
rect 1118 126 1122 130
rect 1061 117 1065 121
rect 1143 126 1147 130
rect 1165 126 1169 130
rect 1185 134 1189 138
rect 1195 126 1199 130
rect 1133 116 1137 120
rect 1219 117 1223 121
rect 1252 126 1256 130
rect 1288 129 1292 133
rect 1251 118 1255 122
rect 1268 121 1272 125
rect 1278 119 1282 123
rect 1241 111 1245 115
rect 1327 127 1331 131
rect 1341 120 1345 124
rect 1310 112 1314 116
rect 999 84 1003 88
rect 396 62 400 66
rect 368 25 373 30
rect 388 14 392 18
rect 498 54 502 59
rect 465 42 469 47
rect 461 25 466 30
rect 554 42 558 46
rect 546 25 551 30
rect 1137 69 1141 73
rect 1122 59 1126 63
rect 1223 68 1227 72
rect 1255 67 1259 71
rect 1147 59 1151 63
rect 1169 59 1173 63
rect 1199 59 1203 63
rect 1282 66 1286 70
rect 1256 59 1260 63
rect 1314 73 1318 77
rect 1345 65 1349 69
rect 1292 56 1296 60
rect 1331 58 1335 62
rect 1189 51 1193 55
rect 312 3 319 10
<< m3contact >>
rect 498 374 502 378
rect 517 353 521 357
<< psubstratepcontact >>
rect 144 441 148 445
rect 231 441 235 445
rect 324 441 328 445
rect 536 443 540 447
rect 629 443 633 447
rect 716 443 720 447
rect 38 302 42 306
rect 116 302 120 306
rect 200 302 204 306
rect 270 302 274 306
rect 367 304 371 308
rect 445 304 449 308
rect 529 304 533 308
rect 599 304 603 308
rect 694 307 698 311
rect 772 307 776 311
rect 856 307 860 311
rect 926 307 930 311
rect 131 292 135 296
rect 159 292 163 296
rect 460 294 464 298
rect 488 294 492 298
rect 787 297 791 301
rect 815 297 819 301
rect 37 156 41 160
rect 115 156 119 160
rect 199 156 203 160
rect 269 156 273 160
rect 366 158 370 162
rect 444 158 448 162
rect 528 158 532 162
rect 598 158 602 162
rect 693 161 697 165
rect 771 161 775 165
rect 855 161 859 165
rect 925 161 929 165
rect 130 146 134 150
rect 158 146 162 150
rect 459 148 463 152
rect 487 148 491 152
rect 786 151 790 155
rect 814 151 818 155
rect 331 8 335 12
rect 424 8 428 12
rect 511 8 515 12
<< nsubstratencontact >>
rect 1172 443 1176 447
rect 1226 443 1230 447
rect 1282 443 1286 447
rect 1336 443 1340 447
rect 144 381 148 385
rect 231 381 235 385
rect 324 381 328 385
rect 536 383 540 387
rect 629 383 633 387
rect 716 383 720 387
rect 38 362 42 366
rect 52 362 56 366
rect 66 362 70 366
rect 149 362 153 366
rect 233 362 237 366
rect 270 362 274 366
rect 284 362 288 366
rect 298 362 302 366
rect 367 364 371 368
rect 381 364 385 368
rect 395 364 399 368
rect 478 364 482 368
rect 562 364 566 368
rect 599 364 603 368
rect 613 364 617 368
rect 627 364 631 368
rect 694 367 698 371
rect 708 367 712 371
rect 722 367 726 371
rect 805 367 809 371
rect 889 367 893 371
rect 926 367 930 371
rect 940 367 944 371
rect 954 367 958 371
rect 1176 316 1180 320
rect 1230 316 1234 320
rect 1286 316 1290 320
rect 1340 316 1344 320
rect 1172 298 1176 302
rect 1226 298 1230 302
rect 1282 298 1286 302
rect 1336 298 1340 302
rect 159 232 163 236
rect 488 234 492 238
rect 815 237 819 241
rect 37 216 41 220
rect 51 216 55 220
rect 65 216 69 220
rect 148 216 152 220
rect 232 216 236 220
rect 269 216 273 220
rect 283 216 287 220
rect 297 216 301 220
rect 366 218 370 222
rect 380 218 384 222
rect 394 218 398 222
rect 477 218 481 222
rect 561 218 565 222
rect 598 218 602 222
rect 612 218 616 222
rect 626 218 630 222
rect 693 221 697 225
rect 707 221 711 225
rect 721 221 725 225
rect 804 221 808 225
rect 888 221 892 225
rect 925 221 929 225
rect 939 221 943 225
rect 953 221 957 225
rect 1176 171 1180 175
rect 1230 171 1234 175
rect 1286 171 1290 175
rect 1340 171 1344 175
rect 1171 156 1175 160
rect 1225 156 1229 160
rect 1281 156 1285 160
rect 1335 156 1339 160
rect 158 86 162 90
rect 487 88 491 92
rect 814 91 818 95
rect 331 68 335 72
rect 424 68 428 72
rect 511 68 515 72
rect 1175 29 1179 33
rect 1229 29 1233 33
rect 1285 29 1289 33
rect 1339 29 1343 33
<< psubstratepdiff >>
rect 535 447 541 448
rect 143 445 149 446
rect 143 441 144 445
rect 148 441 149 445
rect 143 440 149 441
rect 230 445 236 446
rect 230 441 231 445
rect 235 441 236 445
rect 230 440 236 441
rect 323 445 329 446
rect 323 441 324 445
rect 328 441 329 445
rect 535 443 536 447
rect 540 443 541 447
rect 535 442 541 443
rect 628 447 634 448
rect 628 443 629 447
rect 633 443 634 447
rect 323 440 329 441
rect 628 442 634 443
rect 715 447 721 448
rect 715 443 716 447
rect 720 443 721 447
rect 715 442 721 443
rect 37 306 43 307
rect 37 302 38 306
rect 42 302 43 306
rect 37 301 43 302
rect 115 306 121 307
rect 115 302 116 306
rect 120 302 121 306
rect 115 301 121 302
rect 199 306 205 307
rect 199 302 200 306
rect 204 302 205 306
rect 199 301 205 302
rect 366 308 372 309
rect 269 306 275 307
rect 269 302 270 306
rect 274 302 275 306
rect 269 301 275 302
rect 366 304 367 308
rect 371 304 372 308
rect 366 303 372 304
rect 444 308 450 309
rect 444 304 445 308
rect 449 304 450 308
rect 444 303 450 304
rect 528 308 534 309
rect 528 304 529 308
rect 533 304 534 308
rect 528 303 534 304
rect 693 311 699 312
rect 598 308 604 309
rect 598 304 599 308
rect 603 304 604 308
rect 598 303 604 304
rect 693 307 694 311
rect 698 307 699 311
rect 693 306 699 307
rect 771 311 777 312
rect 771 307 772 311
rect 776 307 777 311
rect 771 306 777 307
rect 855 311 861 312
rect 855 307 856 311
rect 860 307 861 311
rect 855 306 861 307
rect 925 311 931 312
rect 925 307 926 311
rect 930 307 931 311
rect 925 306 931 307
rect 786 301 820 302
rect 459 298 493 299
rect 130 296 164 297
rect 130 292 131 296
rect 135 292 159 296
rect 163 292 164 296
rect 459 294 460 298
rect 464 294 488 298
rect 492 294 493 298
rect 786 297 787 301
rect 791 297 815 301
rect 819 297 820 301
rect 786 296 820 297
rect 459 293 493 294
rect 130 291 164 292
rect 36 160 42 161
rect 36 156 37 160
rect 41 156 42 160
rect 36 155 42 156
rect 114 160 120 161
rect 114 156 115 160
rect 119 156 120 160
rect 114 155 120 156
rect 198 160 204 161
rect 198 156 199 160
rect 203 156 204 160
rect 198 155 204 156
rect 365 162 371 163
rect 268 160 274 161
rect 268 156 269 160
rect 273 156 274 160
rect 268 155 274 156
rect 365 158 366 162
rect 370 158 371 162
rect 365 157 371 158
rect 443 162 449 163
rect 443 158 444 162
rect 448 158 449 162
rect 443 157 449 158
rect 527 162 533 163
rect 527 158 528 162
rect 532 158 533 162
rect 527 157 533 158
rect 692 165 698 166
rect 597 162 603 163
rect 597 158 598 162
rect 602 158 603 162
rect 597 157 603 158
rect 692 161 693 165
rect 697 161 698 165
rect 692 160 698 161
rect 770 165 776 166
rect 770 161 771 165
rect 775 161 776 165
rect 770 160 776 161
rect 854 165 860 166
rect 854 161 855 165
rect 859 161 860 165
rect 854 160 860 161
rect 924 165 930 166
rect 924 161 925 165
rect 929 161 930 165
rect 924 160 930 161
rect 785 155 819 156
rect 458 152 492 153
rect 129 150 163 151
rect 129 146 130 150
rect 134 146 158 150
rect 162 146 163 150
rect 458 148 459 152
rect 463 148 487 152
rect 491 148 492 152
rect 785 151 786 155
rect 790 151 814 155
rect 818 151 819 155
rect 785 150 819 151
rect 458 147 492 148
rect 129 145 163 146
rect 330 12 336 13
rect 330 8 331 12
rect 335 8 336 12
rect 330 7 336 8
rect 423 12 429 13
rect 423 8 424 12
rect 428 8 429 12
rect 423 7 429 8
rect 510 12 516 13
rect 510 8 511 12
rect 515 8 516 12
rect 510 7 516 8
<< nsubstratendiff >>
rect 143 385 149 386
rect 230 385 236 386
rect 535 387 541 388
rect 628 387 634 388
rect 715 387 721 388
rect 323 385 329 386
rect 143 381 144 385
rect 148 381 149 385
rect 143 380 149 381
rect 230 381 231 385
rect 235 381 236 385
rect 230 380 236 381
rect 323 381 324 385
rect 328 381 329 385
rect 535 383 536 387
rect 540 383 541 387
rect 535 382 541 383
rect 628 383 629 387
rect 633 383 634 387
rect 628 382 634 383
rect 715 383 716 387
rect 720 383 721 387
rect 715 382 721 383
rect 323 380 329 381
rect 366 368 400 369
rect 37 366 71 367
rect 37 362 38 366
rect 42 362 52 366
rect 56 362 66 366
rect 70 362 71 366
rect 148 366 154 367
rect 37 361 71 362
rect 148 362 149 366
rect 153 362 154 366
rect 232 366 238 367
rect 148 361 154 362
rect 232 362 233 366
rect 237 362 238 366
rect 269 366 303 367
rect 232 361 238 362
rect 269 362 270 366
rect 274 362 284 366
rect 288 362 298 366
rect 302 362 303 366
rect 366 364 367 368
rect 371 364 381 368
rect 385 364 395 368
rect 399 364 400 368
rect 477 368 483 369
rect 366 363 400 364
rect 269 361 303 362
rect 477 364 478 368
rect 482 364 483 368
rect 561 368 567 369
rect 477 363 483 364
rect 561 364 562 368
rect 566 364 567 368
rect 598 368 632 369
rect 561 363 567 364
rect 598 364 599 368
rect 603 364 613 368
rect 617 364 627 368
rect 631 364 632 368
rect 693 367 694 371
rect 698 367 708 371
rect 712 367 722 371
rect 726 367 727 371
rect 804 371 810 372
rect 693 366 727 367
rect 598 363 632 364
rect 804 367 805 371
rect 809 367 810 371
rect 888 371 894 372
rect 804 366 810 367
rect 888 367 889 371
rect 893 367 894 371
rect 925 371 959 372
rect 888 366 894 367
rect 925 367 926 371
rect 930 367 940 371
rect 944 367 954 371
rect 958 367 959 371
rect 925 366 959 367
rect 158 236 164 237
rect 814 241 820 242
rect 487 238 493 239
rect 158 232 159 236
rect 163 232 164 236
rect 487 234 488 238
rect 492 234 493 238
rect 814 237 815 241
rect 819 237 820 241
rect 814 236 820 237
rect 487 233 493 234
rect 158 231 164 232
rect 692 225 726 226
rect 365 222 399 223
rect 36 220 70 221
rect 36 216 37 220
rect 41 216 51 220
rect 55 216 65 220
rect 69 216 70 220
rect 147 220 153 221
rect 36 215 70 216
rect 147 216 148 220
rect 152 216 153 220
rect 231 220 237 221
rect 147 215 153 216
rect 231 216 232 220
rect 236 216 237 220
rect 268 220 302 221
rect 231 215 237 216
rect 268 216 269 220
rect 273 216 283 220
rect 287 216 297 220
rect 301 216 302 220
rect 365 218 366 222
rect 370 218 380 222
rect 384 218 394 222
rect 398 218 399 222
rect 476 222 482 223
rect 365 217 399 218
rect 268 215 302 216
rect 476 218 477 222
rect 481 218 482 222
rect 560 222 566 223
rect 476 217 482 218
rect 560 218 561 222
rect 565 218 566 222
rect 597 222 631 223
rect 560 217 566 218
rect 597 218 598 222
rect 602 218 612 222
rect 616 218 626 222
rect 630 218 631 222
rect 692 221 693 225
rect 697 221 707 225
rect 711 221 721 225
rect 725 221 726 225
rect 803 225 809 226
rect 692 220 726 221
rect 597 217 631 218
rect 803 221 804 225
rect 808 221 809 225
rect 887 225 893 226
rect 803 220 809 221
rect 887 221 888 225
rect 892 221 893 225
rect 924 225 958 226
rect 887 220 893 221
rect 924 221 925 225
rect 929 221 939 225
rect 943 221 953 225
rect 957 221 958 225
rect 924 220 958 221
rect 157 90 163 91
rect 813 95 819 96
rect 486 92 492 93
rect 157 86 158 90
rect 162 86 163 90
rect 486 88 487 92
rect 491 88 492 92
rect 813 91 814 95
rect 818 91 819 95
rect 813 90 819 91
rect 486 87 492 88
rect 157 85 163 86
rect 330 72 336 73
rect 330 68 331 72
rect 335 68 336 72
rect 423 72 429 73
rect 423 68 424 72
rect 428 68 429 72
rect 510 72 516 73
rect 510 68 511 72
rect 515 68 516 72
rect 330 67 336 68
rect 423 67 429 68
rect 510 67 516 68
<< pad >>
rect 171 375 175 379
<< labels >>
rlabel metal1 476 298 476 298 2 vss
rlabel metal1 710 307 710 307 6 vss
rlabel metal1 942 371 942 371 6 vdd
rlabel metal1 803 301 803 301 2 vss
rlabel metal1 803 237 803 237 2 vdd
rlabel metal1 802 91 802 91 2 vdd
rlabel metal1 802 155 802 155 2 vss
rlabel metal1 941 161 941 161 6 vss
rlabel metal1 941 225 941 225 6 vdd
rlabel metal1 709 225 709 225 6 vdd
rlabel metal1 709 161 709 161 6 vss
rlabel metal1 799 225 799 225 6 vdd
rlabel metal1 475 152 475 152 2 vss
rlabel metal1 614 158 614 158 6 vss
rlabel metal1 614 222 614 222 6 vdd
rlabel metal1 382 222 382 222 6 vdd
rlabel metal1 382 158 382 158 6 vss
rlabel metal1 556 222 556 222 6 vdd
rlabel metal1 556 158 556 158 6 vss
rlabel metal1 146 86 146 86 2 vdd
rlabel metal1 53 220 53 220 6 vdd
rlabel metal1 53 156 53 156 6 vss
rlabel metal1 227 220 227 220 6 vdd
rlabel metal1 227 156 227 156 6 vss
rlabel m2contact 112 425 112 425 1 q0_M1
rlabel metal1 148 417 148 417 1 q0b2_M1
rlabel metal1 320 424 320 424 1 q0b0_n_M1
rlabel metal1 440 430 440 430 1 b2_M1
rlabel metal1 441 409 441 409 1 b1_M1
rlabel metal1 441 390 441 390 1 b0_M1
rlabel metal1 535 428 535 428 1 q1b0_M1
rlabel metal1 637 435 637 435 1 q1b1_M1
rlabel metal1 637 413 637 413 1 q1b1_n_M1
rlabel metal1 715 424 715 424 1 q1b2_M1
rlabel metal1 724 424 724 424 1 q1b2_n_M1
rlabel m2contact 751 427 751 427 1 q1_M1
rlabel metal1 940 335 940 335 1 zc1_n_3_M1
rlabel metal1 926 335 926 335 1 c1_3_M1
rlabel metal1 912 339 912 339 1 s_fa3_M1
rlabel metal1 889 357 889 357 1 cn_3_M1
rlabel ntransistor 905 322 905 322 1 s_fa3_n_M1
rlabel metal1 828 339 828 339 1 so_3_M1
rlabel metal1 816 360 816 360 1 bn3_M1
rlabel ptransistor 812 344 812 344 1 an3_M1
rlabel metal1 715 339 715 339 1 co_n3_M1
rlabel metal1 702 319 702 319 1 co_3_M1
rlabel metal1 599 332 599 332 1 c1_2_M1
rlabel metal1 613 332 613 332 1 zc1_2_n_M1
rlabel ntransistor 578 319 578 319 1 son_2_M1
rlabel pdcontact 575 349 575 349 1 s_fa2_M1
rlabel metal1 563 332 563 332 1 cn2_M1
rlabel metal1 501 336 501 336 1 so_2_M1
rlabel polycontact 491 332 491 332 1 an_2_M1
rlabel polycontact 485 333 485 333 1 bn_2_M1
rlabel metal1 388 335 388 335 1 co_n2_M1
rlabel metal1 375 316 375 316 1 co_2_M1
rlabel metal1 284 330 284 330 1 zc1_n1_M1
rlabel metal1 270 330 270 330 1 c1_1_M1
rlabel metal1 256 334 256 334 1 a1_M1
rlabel ntransistor 249 317 249 317 1 a1_n_M1
rlabel ntransistor 165 318 165 318 1 an_1_M1
rlabel metal1 172 334 172 334 1 so_1_M1
rlabel metal1 160 355 160 355 1 bn_1_M1
rlabel metal1 59 334 59 334 1 co_n1_M1
rlabel metal1 46 314 46 314 1 co_1_M1
rlabel metal1 155 262 155 262 1 c_fa1_n_M1
rlabel metal1 163 262 163 262 1 c_fa1_M1
rlabel metal1 484 266 484 266 1 c_fa_n_M1
rlabel metal1 492 270 492 270 1 c_fa2_M1
rlabel metal1 811 269 811 269 1 c_fa3_n_M1
rlabel metal1 819 273 819 273 1 c_fa3_M1
rlabel metal1 939 189 939 189 1 zc1_6_n_M1
rlabel metal1 925 189 925 189 1 c1_6_M1
rlabel ntransistor 904 176 904 176 1 s_fa_6_n_M1
rlabel metal1 911 193 911 193 1 a2_M1
rlabel metal1 887 210 887 210 1 cn_6_M1
rlabel metal1 827 193 827 193 1 so_6_M1
rlabel ptransistor 811 198 811 198 1 an_6_M1
rlabel metal1 772 187 772 187 1 bn_6_M1
rlabel metal1 714 193 714 193 1 co_n_6_M1
rlabel metal1 701 173 701 173 1 co_6_M1
rlabel metal1 612 186 612 186 1 zc1_n_5_M1
rlabel metal1 598 186 598 186 1 c1_5_M1
rlabel metal1 560 206 560 206 1 cn_5_M1
rlabel metal1 584 190 584 190 1 a3_M1
rlabel ntransistor 577 173 577 173 1 s_fa5_n_M1
rlabel metal1 488 211 488 211 1 bn_5_M1
rlabel ptransistor 484 195 484 195 1 an_5_M1
rlabel metal1 500 190 500 190 1 so_5_M1
rlabel metal1 387 190 387 190 1 co_5__M1
rlabel metal1 283 184 283 184 1 zc1_4_M1
rlabel metal1 269 184 269 184 1 c1_4_M1
rlabel metal1 255 188 255 188 1 a4_M1
rlabel ntransistor 248 171 248 171 1 s_fa4_n_M1
rlabel metal1 231 204 231 204 1 cn_1_M1
rlabel metal1 148 203 148 203 1 bn4_M1
rlabel ptransistor 155 193 155 193 1 an4_M1
rlabel metal1 171 188 171 188 1 so_4_M1
rlabel metal1 58 188 58 188 1 co_n4_M1
rlabel metal1 45 168 45 168 1 co_4_M1
rlabel metal1 154 118 154 118 1 a5_n_M1
rlabel metal1 162 122 162 122 1 a5_M1
rlabel metal1 491 124 491 124 1 c_fa5_M1
rlabel metal1 483 120 483 120 1 c_fa5_n_M1
rlabel metal1 810 123 810 123 1 c_fa6_n_M1
rlabel metal1 818 127 818 127 1 c_fa6_M1
rlabel metal1 511 30 511 30 1 q2b0_M1
rlabel metal1 520 29 520 29 1 q2b0_n_M1
rlabel m2contact 548 28 548 28 1 q2_M1
rlabel metal1 423 30 423 30 1 q2b1_M1
rlabel metal1 432 30 432 30 1 q2b1_n_M1
rlabel metal1 353 19 353 19 1 q2b2_n_M1
rlabel metal1 331 18 331 18 1 q2b2_M1
rlabel metal1 140 421 140 421 1 q0b2_n_M1
rlabel metal1 235 421 235 421 1 q0b1_M1
rlabel metal1 544 414 544 414 1 q1b0_n_M1
rlabel metal1 227 422 227 422 1 q0b1_n_M1
rlabel metal1 327 423 327 423 1 a0_M1
rlabel metal1 1332 310 1332 310 1 vdd
rlabel m2contact 1063 406 1063 406 1 en_bar_D1
rlabel metal1 1134 413 1134 413 1 D_bar_D1
rlabel polycontact 1173 414 1173 414 1 en_D1
rlabel metal1 1181 411 1181 411 1 out_n1_D1
rlabel ndiffusion 1162 394 1162 394 1 n1_D1
rlabel ndiffusion 1218 394 1218 394 1 n2_D1
rlabel metal1 1236 407 1236 407 1 out_n2_D1
rlabel ndiffusion 1274 394 1274 394 1 n3_D1
rlabel ndiffusion 1328 394 1328 394 1 n4_D1
rlabel m2contact 1345 410 1345 410 1 q_l1_bar_D1
rlabel m2contact 1349 353 1349 353 1 q_bar_D1
rlabel ndiffusion 1332 369 1332 369 1 n10_D1
rlabel metal1 1240 356 1240 356 1 out_n8_D1
rlabel ndiffusion 1222 369 1222 369 1 n8_D1
rlabel metal1 1185 352 1185 352 1 out_n7_D1
rlabel ndiffusion 1166 369 1166 369 1 n7_D1
rlabel polycontact 1156 349 1156 349 1 q_l1_D1
rlabel metal1 1138 353 1138 353 1 n6_D1
rlabel ndiffusion 1278 369 1278 369 1 n9_D1
rlabel m2contact 1295 345 1295 345 1 q_D1
rlabel metal2 1398 306 1398 306 8 q_D1
rlabel m2contact 1345 265 1345 265 1 q_l1_bar_D2
rlabel metal1 1138 208 1138 208 1 n6_D2
rlabel polycontact 1156 204 1156 204 1 q_l1_D2
rlabel ndiffusion 1166 224 1166 224 1 n7_D2
rlabel metal1 1185 207 1185 207 1 out_n7__D2
rlabel ndiffusion 1222 224 1222 224 1 n8_D2
rlabel metal1 1240 211 1240 211 1 out_n8_D2
rlabel ndiffusion 1278 224 1278 224 1 n9_D2
rlabel m2contact 1295 200 1295 200 1 q_D2
rlabel ndiffusion 1332 224 1332 224 1 n10_D2
rlabel m2contact 1349 208 1349 208 1 q_bar_D2
rlabel ndiffusion 1328 249 1328 249 1 n4_D2
rlabel ndiffusion 1274 249 1274 249 1 n3_D2
rlabel metal1 1236 262 1236 262 1 out_n2_D2
rlabel ndiffusion 1218 249 1218 249 1 n2_D2
rlabel metal1 1181 266 1181 266 1 out_n1_D2
rlabel ndiffusion 1162 249 1162 249 1 n1_D2
rlabel metal1 1134 268 1134 268 1 D_bar_D2
rlabel m2contact 1063 261 1063 261 1 en_bar_D2
rlabel metal1 1332 165 1332 165 1 vdd
rlabel metal1 1172 97 1172 97 1 vss
rlabel metal1 1137 66 1137 66 1 n6_D3
rlabel polycontact 1155 62 1155 62 1 q_l1_D3
rlabel ndiffusion 1165 82 1165 82 1 n7_D3
rlabel metal1 1184 65 1184 65 1 out_n7_D3
rlabel ndiffusion 1221 82 1221 82 1 n8_D3
rlabel m2contact 1294 58 1294 58 1 q_D3
rlabel metal1 1239 69 1239 69 1 out_n8_D3
rlabel ndiffusion 1277 82 1277 82 1 n9_D3
rlabel m2contact 1348 66 1348 66 1 q_bar_D3
rlabel m2contact 1344 123 1344 123 1 q_l1_bar_D3
rlabel ndiffusion 1327 107 1327 107 1 n4_D3
rlabel ndiffusion 1273 107 1273 107 1 n3_D3
rlabel metal1 1235 120 1235 120 1 out_n2_D3
rlabel ndiffusion 1217 107 1217 107 1 n2_D3
rlabel metal1 1180 124 1180 124 1 out_n1_D3
rlabel ndiffusion 1161 107 1161 107 1 n1_D3
rlabel metal1 1133 126 1133 126 1 D_bar_D3
rlabel m2contact 1062 119 1062 119 1 en_bar_D3
rlabel ndiffusion 1331 82 1331 82 1 n10
rlabel metal1 1331 23 1331 23 1 vdd
rlabel metal2 1369 172 1369 172 1 q_D2
rlabel metal2 1367 27 1367 27 1 q_D3
<< end >>
