magic
tech scmos
timestamp 1523024729
<< pwell >>
rect -708 -72 -690 -68
rect -710 -76 -690 -72
rect -710 -112 -662 -76
rect -623 -112 -575 -76
rect -530 -112 -482 -76
rect -290 -110 -242 -74
rect -197 -110 -149 -74
rect -110 -110 -62 -74
rect -781 -235 -638 -199
rect -626 -235 -508 -199
rect -452 -233 -309 -197
rect -297 -233 -179 -197
rect -125 -230 18 -194
rect 30 -230 148 -194
rect -695 -261 -647 -235
rect -366 -259 -318 -233
rect -39 -256 9 -230
rect -782 -381 -639 -345
rect -627 -381 -509 -345
rect -453 -379 -310 -343
rect -298 -379 -180 -343
rect -126 -376 17 -340
rect 29 -376 147 -340
rect -696 -407 -648 -381
rect -367 -405 -319 -379
rect -40 -402 8 -376
rect -495 -529 -447 -493
rect -402 -529 -354 -493
rect -315 -529 -267 -493
<< nwell >>
rect -115 -42 64 -16
rect 77 -42 118 -16
rect 133 -42 174 -16
rect 187 -42 228 -16
rect -710 -155 -662 -112
rect -623 -155 -575 -112
rect -530 -155 -482 -112
rect -290 -147 -242 -110
rect -197 -147 -149 -110
rect -290 -150 -149 -147
rect -294 -153 -149 -150
rect -110 -141 -62 -110
rect -19 -140 68 -121
rect 81 -140 122 -121
rect 137 -140 178 -121
rect -110 -150 -49 -141
rect -25 -147 178 -140
rect 191 -147 232 -121
rect -25 -149 160 -147
rect -25 -150 157 -149
rect -110 -153 157 -150
rect -781 -199 -638 -155
rect -626 -156 -482 -155
rect -626 -199 -508 -156
rect -452 -197 -309 -153
rect -297 -157 157 -153
rect -297 -167 18 -157
rect -297 -197 -179 -167
rect -125 -194 18 -167
rect 30 -159 157 -157
rect 30 -194 148 -159
rect -695 -268 -647 -261
rect -366 -266 -318 -259
rect -39 -263 9 -256
rect -699 -281 -647 -268
rect -370 -279 -318 -266
rect -43 -276 9 -263
rect -695 -297 -647 -281
rect -366 -295 -318 -279
rect -39 -289 9 -276
rect -706 -301 -640 -297
rect -376 -299 -310 -295
rect -68 -296 43 -289
rect -782 -345 -639 -301
rect -627 -345 -509 -301
rect -453 -343 -310 -299
rect -298 -343 -180 -299
rect -126 -305 147 -296
rect -126 -340 17 -305
rect 29 -340 147 -305
rect -696 -414 -648 -407
rect -367 -412 -319 -405
rect -40 -409 8 -402
rect -700 -427 -648 -414
rect -371 -425 -319 -412
rect -44 -422 8 -409
rect -696 -451 -648 -427
rect -367 -435 -319 -425
rect -493 -449 -261 -435
rect -40 -446 8 -422
rect -495 -452 -261 -449
rect -495 -493 -447 -452
rect -402 -493 -354 -452
rect -315 -493 -267 -452
<< polysilicon >>
rect -78 -29 -76 -27
rect -6 -29 -4 -23
rect 33 -29 35 -23
rect 54 -29 56 -23
rect 87 -29 89 -23
rect 108 -29 110 -23
rect 143 -29 145 -23
rect 164 -29 166 -23
rect 197 -29 199 -23
rect 218 -29 220 -23
rect -78 -46 -76 -35
rect -6 -47 -4 -35
rect 33 -47 35 -35
rect 54 -47 56 -35
rect 87 -47 89 -35
rect 108 -47 110 -35
rect 143 -47 145 -35
rect 164 -47 166 -35
rect 197 -47 199 -35
rect 218 -47 220 -35
rect -78 -68 -76 -50
rect 34 -51 35 -47
rect 55 -51 56 -47
rect 88 -51 89 -47
rect 109 -51 110 -47
rect 144 -51 145 -47
rect 165 -51 166 -47
rect 198 -51 199 -47
rect 219 -51 220 -47
rect -78 -74 -76 -71
rect -6 -69 -4 -51
rect 33 -66 35 -51
rect 54 -66 56 -51
rect 87 -66 89 -51
rect 108 -66 110 -51
rect 143 -66 145 -51
rect 164 -66 166 -51
rect 197 -66 199 -51
rect 218 -66 220 -51
rect -6 -75 -4 -72
rect 33 -75 35 -72
rect 54 -75 56 -72
rect 87 -75 89 -72
rect 108 -75 110 -72
rect 143 -75 145 -72
rect 164 -75 166 -72
rect 197 -75 199 -72
rect 218 -75 220 -72
rect -697 -93 -695 -88
rect -690 -93 -688 -88
rect -677 -95 -675 -91
rect -610 -93 -608 -88
rect -603 -93 -601 -88
rect -590 -95 -588 -91
rect -517 -93 -515 -88
rect -510 -93 -508 -88
rect -497 -95 -495 -91
rect -277 -93 -275 -89
rect -264 -91 -262 -86
rect -257 -91 -255 -86
rect -184 -93 -182 -89
rect -171 -91 -169 -86
rect -164 -91 -162 -86
rect -97 -93 -95 -89
rect -84 -91 -82 -86
rect -77 -91 -75 -86
rect -2 -91 0 -88
rect 37 -91 39 -88
rect 58 -91 60 -88
rect 91 -91 93 -88
rect 112 -91 114 -88
rect 147 -91 149 -88
rect 168 -91 170 -88
rect 201 -91 203 -88
rect 222 -91 224 -88
rect -697 -117 -695 -104
rect -690 -109 -688 -104
rect -677 -109 -675 -104
rect -691 -110 -685 -109
rect -691 -114 -690 -110
rect -686 -114 -685 -110
rect -691 -115 -685 -114
rect -681 -110 -675 -109
rect -681 -114 -680 -110
rect -676 -114 -675 -110
rect -681 -115 -675 -114
rect -701 -118 -695 -117
rect -701 -122 -700 -118
rect -696 -122 -695 -118
rect -701 -123 -695 -122
rect -697 -126 -695 -123
rect -687 -126 -685 -115
rect -677 -119 -675 -115
rect -610 -117 -608 -104
rect -603 -109 -601 -104
rect -590 -109 -588 -104
rect -604 -110 -598 -109
rect -604 -114 -603 -110
rect -599 -114 -598 -110
rect -604 -115 -598 -114
rect -594 -110 -588 -109
rect -594 -114 -593 -110
rect -589 -114 -588 -110
rect -594 -115 -588 -114
rect -614 -118 -608 -117
rect -614 -122 -613 -118
rect -609 -122 -608 -118
rect -614 -123 -608 -122
rect -610 -126 -608 -123
rect -600 -126 -598 -115
rect -590 -119 -588 -115
rect -517 -117 -515 -104
rect -510 -109 -508 -104
rect -497 -109 -495 -104
rect -511 -110 -505 -109
rect -511 -114 -510 -110
rect -506 -114 -505 -110
rect -511 -115 -505 -114
rect -501 -110 -495 -109
rect -501 -114 -500 -110
rect -496 -114 -495 -110
rect -501 -115 -495 -114
rect -521 -118 -515 -117
rect -697 -144 -695 -139
rect -687 -144 -685 -139
rect -677 -141 -675 -137
rect -521 -122 -520 -118
rect -516 -122 -515 -118
rect -521 -123 -515 -122
rect -517 -126 -515 -123
rect -507 -126 -505 -115
rect -497 -119 -495 -115
rect -277 -107 -275 -102
rect -264 -107 -262 -102
rect -277 -108 -271 -107
rect -277 -112 -276 -108
rect -272 -112 -271 -108
rect -277 -113 -271 -112
rect -267 -108 -261 -107
rect -267 -112 -266 -108
rect -262 -112 -261 -108
rect -267 -113 -261 -112
rect -277 -117 -275 -113
rect -610 -144 -608 -139
rect -600 -144 -598 -139
rect -590 -141 -588 -137
rect -267 -124 -265 -113
rect -257 -115 -255 -102
rect -184 -107 -182 -102
rect -171 -107 -169 -102
rect -184 -108 -178 -107
rect -184 -112 -183 -108
rect -179 -112 -178 -108
rect -184 -113 -178 -112
rect -174 -108 -168 -107
rect -174 -112 -173 -108
rect -169 -112 -168 -108
rect -174 -113 -168 -112
rect -257 -116 -251 -115
rect -257 -120 -256 -116
rect -252 -120 -251 -116
rect -184 -117 -182 -113
rect -257 -121 -251 -120
rect -257 -124 -255 -121
rect -517 -144 -515 -139
rect -507 -144 -505 -139
rect -497 -141 -495 -137
rect -277 -139 -275 -135
rect -174 -124 -172 -113
rect -164 -115 -162 -102
rect -97 -107 -95 -102
rect -84 -107 -82 -102
rect -97 -108 -91 -107
rect -97 -112 -96 -108
rect -92 -112 -91 -108
rect -97 -113 -91 -112
rect -87 -108 -81 -107
rect -87 -112 -86 -108
rect -82 -112 -81 -108
rect -87 -113 -81 -112
rect -164 -116 -158 -115
rect -164 -120 -163 -116
rect -159 -120 -158 -116
rect -97 -117 -95 -113
rect -164 -121 -158 -120
rect -164 -124 -162 -121
rect -267 -142 -265 -137
rect -257 -142 -255 -137
rect -184 -139 -182 -135
rect -87 -124 -85 -113
rect -77 -115 -75 -102
rect -2 -112 0 -94
rect 37 -112 39 -97
rect 58 -112 60 -97
rect 91 -112 93 -97
rect 112 -112 114 -97
rect 147 -112 149 -97
rect 168 -112 170 -97
rect 201 -112 203 -97
rect 222 -112 224 -97
rect -77 -116 -71 -115
rect 38 -116 39 -112
rect 59 -116 60 -112
rect 92 -116 93 -112
rect 113 -116 114 -112
rect 148 -116 149 -112
rect 169 -116 170 -112
rect 202 -116 203 -112
rect 223 -116 224 -112
rect -77 -120 -76 -116
rect -72 -120 -71 -116
rect -77 -121 -71 -120
rect -77 -124 -75 -121
rect -174 -142 -172 -137
rect -164 -142 -162 -137
rect -97 -139 -95 -135
rect -2 -128 0 -116
rect 37 -123 39 -116
rect 37 -128 39 -126
rect 58 -128 60 -116
rect 91 -128 93 -116
rect 112 -128 114 -116
rect 147 -128 149 -116
rect 168 -128 170 -116
rect 201 -128 203 -116
rect 222 -128 224 -116
rect -87 -142 -85 -137
rect -77 -142 -75 -137
rect -2 -140 0 -134
rect 37 -140 39 -134
rect 58 -140 60 -134
rect 91 -140 93 -134
rect 112 -140 114 -134
rect 147 -140 149 -134
rect 168 -140 170 -134
rect 201 -140 203 -134
rect 222 -140 224 -134
rect -689 -165 -687 -161
rect -765 -173 -759 -172
rect -775 -181 -773 -176
rect -765 -177 -764 -173
rect -760 -177 -759 -173
rect -765 -178 -759 -177
rect -765 -183 -763 -178
rect -755 -183 -753 -178
rect -704 -181 -698 -180
rect -704 -185 -703 -181
rect -699 -185 -698 -181
rect -704 -186 -698 -185
rect -775 -196 -773 -193
rect -765 -196 -763 -193
rect -775 -197 -769 -196
rect -775 -201 -774 -197
rect -770 -201 -769 -197
rect -765 -199 -761 -196
rect -775 -202 -769 -201
rect -775 -210 -773 -202
rect -763 -213 -761 -199
rect -755 -204 -753 -193
rect -700 -195 -698 -186
rect -653 -165 -651 -161
rect -605 -165 -603 -161
rect -673 -174 -671 -170
rect -663 -174 -661 -170
rect -620 -181 -614 -180
rect -620 -185 -619 -181
rect -615 -185 -614 -181
rect -620 -186 -614 -185
rect -689 -195 -687 -192
rect -673 -195 -671 -192
rect -663 -195 -661 -192
rect -653 -195 -651 -192
rect -700 -197 -687 -195
rect -681 -197 -671 -195
rect -667 -196 -661 -195
rect -756 -205 -750 -204
rect -697 -205 -695 -197
rect -681 -201 -679 -197
rect -667 -200 -666 -196
rect -662 -200 -661 -196
rect -667 -201 -661 -200
rect -657 -196 -651 -195
rect -657 -200 -656 -196
rect -652 -200 -651 -196
rect -616 -195 -614 -186
rect -569 -165 -567 -161
rect -589 -174 -587 -170
rect -579 -174 -577 -170
rect -360 -163 -358 -159
rect -436 -171 -430 -170
rect -533 -173 -527 -172
rect -543 -181 -541 -176
rect -533 -177 -532 -173
rect -528 -177 -527 -173
rect -533 -178 -527 -177
rect -605 -195 -603 -192
rect -589 -195 -587 -192
rect -579 -195 -577 -192
rect -569 -195 -567 -192
rect -533 -183 -531 -178
rect -523 -183 -521 -178
rect -446 -179 -444 -174
rect -436 -175 -435 -171
rect -431 -175 -430 -171
rect -436 -176 -430 -175
rect -436 -181 -434 -176
rect -426 -181 -424 -176
rect -375 -179 -369 -178
rect -375 -183 -374 -179
rect -370 -183 -369 -179
rect -375 -184 -369 -183
rect -616 -197 -603 -195
rect -597 -197 -587 -195
rect -583 -196 -577 -195
rect -657 -201 -651 -200
rect -688 -202 -679 -201
rect -756 -209 -755 -205
rect -751 -209 -750 -205
rect -756 -210 -750 -209
rect -756 -213 -754 -210
rect -775 -220 -773 -216
rect -688 -206 -687 -202
rect -683 -206 -679 -202
rect -663 -205 -661 -201
rect -688 -207 -679 -206
rect -681 -210 -679 -207
rect -671 -210 -669 -205
rect -663 -207 -659 -205
rect -661 -210 -659 -207
rect -654 -210 -652 -201
rect -613 -205 -611 -197
rect -597 -201 -595 -197
rect -583 -200 -582 -196
rect -578 -200 -577 -196
rect -583 -201 -577 -200
rect -573 -196 -567 -195
rect -573 -200 -572 -196
rect -568 -200 -567 -196
rect -573 -201 -567 -200
rect -543 -196 -541 -193
rect -533 -196 -531 -193
rect -543 -197 -537 -196
rect -543 -201 -542 -197
rect -538 -201 -537 -197
rect -533 -199 -529 -196
rect -604 -202 -595 -201
rect -697 -217 -695 -214
rect -697 -219 -692 -217
rect -763 -227 -761 -222
rect -756 -227 -754 -222
rect -694 -227 -692 -219
rect -681 -223 -679 -219
rect -671 -227 -669 -219
rect -604 -206 -603 -202
rect -599 -206 -595 -202
rect -579 -205 -577 -201
rect -604 -207 -595 -206
rect -597 -210 -595 -207
rect -587 -210 -585 -205
rect -579 -207 -575 -205
rect -577 -210 -575 -207
rect -570 -210 -568 -201
rect -543 -202 -537 -201
rect -543 -210 -541 -202
rect -613 -217 -611 -214
rect -613 -219 -608 -217
rect -661 -227 -659 -222
rect -654 -227 -652 -222
rect -694 -229 -669 -227
rect -610 -227 -608 -219
rect -597 -223 -595 -219
rect -587 -227 -585 -219
rect -531 -213 -529 -199
rect -523 -204 -521 -193
rect -446 -194 -444 -191
rect -436 -194 -434 -191
rect -446 -195 -440 -194
rect -446 -199 -445 -195
rect -441 -199 -440 -195
rect -436 -197 -432 -194
rect -446 -200 -440 -199
rect -524 -205 -518 -204
rect -524 -209 -523 -205
rect -519 -209 -518 -205
rect -446 -208 -444 -200
rect -524 -210 -518 -209
rect -524 -213 -522 -210
rect -543 -220 -541 -216
rect -434 -211 -432 -197
rect -426 -202 -424 -191
rect -371 -193 -369 -184
rect -324 -163 -322 -159
rect -276 -163 -274 -159
rect -344 -172 -342 -168
rect -334 -172 -332 -168
rect -291 -179 -285 -178
rect -291 -183 -290 -179
rect -286 -183 -285 -179
rect -291 -184 -285 -183
rect -360 -193 -358 -190
rect -344 -193 -342 -190
rect -334 -193 -332 -190
rect -324 -193 -322 -190
rect -371 -195 -358 -193
rect -352 -195 -342 -193
rect -338 -194 -332 -193
rect -427 -203 -421 -202
rect -368 -203 -366 -195
rect -352 -199 -350 -195
rect -338 -198 -337 -194
rect -333 -198 -332 -194
rect -338 -199 -332 -198
rect -328 -194 -322 -193
rect -328 -198 -327 -194
rect -323 -198 -322 -194
rect -287 -193 -285 -184
rect -240 -163 -238 -159
rect -260 -172 -258 -168
rect -250 -172 -248 -168
rect -33 -160 -31 -156
rect -109 -168 -103 -167
rect -204 -171 -198 -170
rect -214 -179 -212 -174
rect -204 -175 -203 -171
rect -199 -175 -198 -171
rect -204 -176 -198 -175
rect -119 -176 -117 -171
rect -109 -172 -108 -168
rect -104 -172 -103 -168
rect -109 -173 -103 -172
rect -276 -193 -274 -190
rect -260 -193 -258 -190
rect -250 -193 -248 -190
rect -240 -193 -238 -190
rect -204 -181 -202 -176
rect -194 -181 -192 -176
rect -109 -178 -107 -173
rect -99 -178 -97 -173
rect -48 -176 -42 -175
rect -48 -180 -47 -176
rect -43 -180 -42 -176
rect -48 -181 -42 -180
rect -119 -191 -117 -188
rect -109 -191 -107 -188
rect -287 -195 -274 -193
rect -268 -195 -258 -193
rect -254 -194 -248 -193
rect -328 -199 -322 -198
rect -359 -200 -350 -199
rect -427 -207 -426 -203
rect -422 -207 -421 -203
rect -427 -208 -421 -207
rect -427 -211 -425 -208
rect -446 -218 -444 -214
rect -359 -204 -358 -200
rect -354 -204 -350 -200
rect -334 -203 -332 -199
rect -359 -205 -350 -204
rect -352 -208 -350 -205
rect -342 -208 -340 -203
rect -334 -205 -330 -203
rect -332 -208 -330 -205
rect -325 -208 -323 -199
rect -284 -203 -282 -195
rect -268 -199 -266 -195
rect -254 -198 -253 -194
rect -249 -198 -248 -194
rect -254 -199 -248 -198
rect -244 -194 -238 -193
rect -244 -198 -243 -194
rect -239 -198 -238 -194
rect -244 -199 -238 -198
rect -214 -194 -212 -191
rect -204 -194 -202 -191
rect -214 -195 -208 -194
rect -214 -199 -213 -195
rect -209 -199 -208 -195
rect -204 -197 -200 -194
rect -275 -200 -266 -199
rect -368 -215 -366 -212
rect -368 -217 -363 -215
rect -577 -227 -575 -222
rect -570 -227 -568 -222
rect -610 -229 -585 -227
rect -531 -227 -529 -222
rect -524 -227 -522 -222
rect -434 -225 -432 -220
rect -427 -225 -425 -220
rect -365 -225 -363 -217
rect -352 -221 -350 -217
rect -342 -225 -340 -217
rect -275 -204 -274 -200
rect -270 -204 -266 -200
rect -250 -203 -248 -199
rect -275 -205 -266 -204
rect -268 -208 -266 -205
rect -258 -208 -256 -203
rect -250 -205 -246 -203
rect -248 -208 -246 -205
rect -241 -208 -239 -199
rect -214 -200 -208 -199
rect -214 -208 -212 -200
rect -284 -215 -282 -212
rect -284 -217 -279 -215
rect -332 -225 -330 -220
rect -325 -225 -323 -220
rect -365 -227 -340 -225
rect -281 -225 -279 -217
rect -268 -221 -266 -217
rect -258 -225 -256 -217
rect -202 -211 -200 -197
rect -194 -202 -192 -191
rect -119 -192 -113 -191
rect -119 -196 -118 -192
rect -114 -196 -113 -192
rect -109 -194 -105 -191
rect -119 -197 -113 -196
rect -195 -203 -189 -202
rect -195 -207 -194 -203
rect -190 -207 -189 -203
rect -119 -205 -117 -197
rect -195 -208 -189 -207
rect -195 -211 -193 -208
rect -107 -208 -105 -194
rect -99 -199 -97 -188
rect -44 -190 -42 -181
rect 3 -160 5 -156
rect 51 -160 53 -156
rect -17 -169 -15 -165
rect -7 -169 -5 -165
rect 36 -176 42 -175
rect 36 -180 37 -176
rect 41 -180 42 -176
rect 36 -181 42 -180
rect -33 -190 -31 -187
rect -17 -190 -15 -187
rect -7 -190 -5 -187
rect 3 -190 5 -187
rect -44 -192 -31 -190
rect -25 -192 -15 -190
rect -11 -191 -5 -190
rect -100 -200 -94 -199
rect -41 -200 -39 -192
rect -25 -196 -23 -192
rect -11 -195 -10 -191
rect -6 -195 -5 -191
rect -11 -196 -5 -195
rect -1 -191 5 -190
rect -1 -195 0 -191
rect 4 -195 5 -191
rect 40 -190 42 -181
rect 87 -160 89 -156
rect 67 -169 69 -165
rect 77 -169 79 -165
rect 123 -168 129 -167
rect 113 -176 115 -171
rect 123 -172 124 -168
rect 128 -172 129 -168
rect 123 -173 129 -172
rect 51 -190 53 -187
rect 67 -190 69 -187
rect 77 -190 79 -187
rect 87 -190 89 -187
rect 123 -178 125 -173
rect 133 -178 135 -173
rect 40 -192 53 -190
rect 59 -192 69 -190
rect 73 -191 79 -190
rect -1 -196 5 -195
rect -32 -197 -23 -196
rect -100 -204 -99 -200
rect -95 -204 -94 -200
rect -100 -205 -94 -204
rect -100 -208 -98 -205
rect -214 -218 -212 -214
rect -119 -215 -117 -211
rect -32 -201 -31 -197
rect -27 -201 -23 -197
rect -7 -200 -5 -196
rect -32 -202 -23 -201
rect -25 -205 -23 -202
rect -15 -205 -13 -200
rect -7 -202 -3 -200
rect -5 -205 -3 -202
rect 2 -205 4 -196
rect 43 -200 45 -192
rect 59 -196 61 -192
rect 73 -195 74 -191
rect 78 -195 79 -191
rect 73 -196 79 -195
rect 83 -191 89 -190
rect 83 -195 84 -191
rect 88 -195 89 -191
rect 83 -196 89 -195
rect 113 -191 115 -188
rect 123 -191 125 -188
rect 113 -192 119 -191
rect 113 -196 114 -192
rect 118 -196 119 -192
rect 123 -194 127 -191
rect 52 -197 61 -196
rect -41 -212 -39 -209
rect -41 -214 -36 -212
rect -248 -225 -246 -220
rect -241 -225 -239 -220
rect -281 -227 -256 -225
rect -202 -225 -200 -220
rect -195 -225 -193 -220
rect -107 -222 -105 -217
rect -100 -222 -98 -217
rect -38 -222 -36 -214
rect -25 -218 -23 -214
rect -15 -222 -13 -214
rect 52 -201 53 -197
rect 57 -201 61 -197
rect 77 -200 79 -196
rect 52 -202 61 -201
rect 59 -205 61 -202
rect 69 -205 71 -200
rect 77 -202 81 -200
rect 79 -205 81 -202
rect 86 -205 88 -196
rect 113 -197 119 -196
rect 113 -205 115 -197
rect 43 -212 45 -209
rect 43 -214 48 -212
rect -5 -222 -3 -217
rect 2 -222 4 -217
rect -38 -224 -13 -222
rect 46 -222 48 -214
rect 59 -218 61 -214
rect 69 -222 71 -214
rect 125 -208 127 -194
rect 133 -199 135 -188
rect 132 -200 138 -199
rect 132 -204 133 -200
rect 137 -204 138 -200
rect 132 -205 138 -204
rect 132 -208 134 -205
rect 113 -215 115 -211
rect 79 -222 81 -217
rect 86 -222 88 -217
rect 46 -224 71 -222
rect 125 -222 127 -217
rect 132 -222 134 -217
rect -682 -244 -680 -240
rect -672 -244 -670 -240
rect -662 -244 -660 -240
rect -353 -242 -351 -238
rect -343 -242 -341 -238
rect -333 -242 -331 -238
rect -26 -239 -24 -235
rect -16 -239 -14 -235
rect -6 -239 -4 -235
rect -682 -258 -680 -250
rect -686 -259 -680 -258
rect -672 -259 -670 -250
rect -662 -259 -660 -250
rect -353 -256 -351 -248
rect -686 -263 -685 -259
rect -681 -263 -680 -259
rect -666 -260 -660 -259
rect -686 -264 -680 -263
rect -682 -277 -680 -264
rect -672 -266 -670 -263
rect -666 -264 -665 -260
rect -661 -264 -660 -260
rect -357 -257 -351 -256
rect -343 -257 -341 -248
rect -333 -257 -331 -248
rect -26 -253 -24 -245
rect -357 -261 -356 -257
rect -352 -261 -351 -257
rect -337 -258 -331 -257
rect -357 -262 -351 -261
rect -666 -265 -660 -264
rect -676 -267 -670 -266
rect -676 -271 -675 -267
rect -671 -271 -670 -267
rect -676 -272 -670 -271
rect -675 -277 -673 -272
rect -662 -274 -660 -265
rect -353 -275 -351 -262
rect -343 -264 -341 -261
rect -337 -262 -336 -258
rect -332 -262 -331 -258
rect -30 -254 -24 -253
rect -16 -254 -14 -245
rect -6 -254 -4 -245
rect -30 -258 -29 -254
rect -25 -258 -24 -254
rect -10 -255 -4 -254
rect -30 -259 -24 -258
rect -337 -263 -331 -262
rect -347 -265 -341 -264
rect -347 -269 -346 -265
rect -342 -269 -341 -265
rect -347 -270 -341 -269
rect -346 -275 -344 -270
rect -333 -272 -331 -263
rect -26 -272 -24 -259
rect -16 -261 -14 -258
rect -10 -259 -9 -255
rect -5 -259 -4 -255
rect -10 -260 -4 -259
rect -20 -262 -14 -261
rect -20 -266 -19 -262
rect -15 -266 -14 -262
rect -20 -267 -14 -266
rect -19 -272 -17 -267
rect -6 -269 -4 -260
rect -662 -290 -660 -286
rect -333 -288 -331 -284
rect -6 -285 -4 -281
rect -682 -299 -680 -295
rect -675 -299 -673 -295
rect -353 -297 -351 -293
rect -346 -297 -344 -293
rect -26 -294 -24 -290
rect -19 -294 -17 -290
rect -690 -311 -688 -307
rect -766 -319 -760 -318
rect -776 -327 -774 -322
rect -766 -323 -765 -319
rect -761 -323 -760 -319
rect -766 -324 -760 -323
rect -766 -329 -764 -324
rect -756 -329 -754 -324
rect -705 -327 -699 -326
rect -705 -331 -704 -327
rect -700 -331 -699 -327
rect -705 -332 -699 -331
rect -776 -342 -774 -339
rect -766 -342 -764 -339
rect -776 -343 -770 -342
rect -776 -347 -775 -343
rect -771 -347 -770 -343
rect -766 -345 -762 -342
rect -776 -348 -770 -347
rect -776 -356 -774 -348
rect -764 -359 -762 -345
rect -756 -350 -754 -339
rect -701 -341 -699 -332
rect -654 -311 -652 -307
rect -606 -311 -604 -307
rect -674 -320 -672 -316
rect -664 -320 -662 -316
rect -621 -327 -615 -326
rect -621 -331 -620 -327
rect -616 -331 -615 -327
rect -621 -332 -615 -331
rect -690 -341 -688 -338
rect -674 -341 -672 -338
rect -664 -341 -662 -338
rect -654 -341 -652 -338
rect -701 -343 -688 -341
rect -682 -343 -672 -341
rect -668 -342 -662 -341
rect -757 -351 -751 -350
rect -698 -351 -696 -343
rect -682 -347 -680 -343
rect -668 -346 -667 -342
rect -663 -346 -662 -342
rect -668 -347 -662 -346
rect -658 -342 -652 -341
rect -658 -346 -657 -342
rect -653 -346 -652 -342
rect -617 -341 -615 -332
rect -570 -311 -568 -307
rect -590 -320 -588 -316
rect -580 -320 -578 -316
rect -361 -309 -359 -305
rect -437 -317 -431 -316
rect -534 -319 -528 -318
rect -544 -327 -542 -322
rect -534 -323 -533 -319
rect -529 -323 -528 -319
rect -534 -324 -528 -323
rect -606 -341 -604 -338
rect -590 -341 -588 -338
rect -580 -341 -578 -338
rect -570 -341 -568 -338
rect -534 -329 -532 -324
rect -524 -329 -522 -324
rect -447 -325 -445 -320
rect -437 -321 -436 -317
rect -432 -321 -431 -317
rect -437 -322 -431 -321
rect -437 -327 -435 -322
rect -427 -327 -425 -322
rect -376 -325 -370 -324
rect -376 -329 -375 -325
rect -371 -329 -370 -325
rect -376 -330 -370 -329
rect -617 -343 -604 -341
rect -598 -343 -588 -341
rect -584 -342 -578 -341
rect -658 -347 -652 -346
rect -689 -348 -680 -347
rect -757 -355 -756 -351
rect -752 -355 -751 -351
rect -757 -356 -751 -355
rect -757 -359 -755 -356
rect -776 -366 -774 -362
rect -689 -352 -688 -348
rect -684 -352 -680 -348
rect -664 -351 -662 -347
rect -689 -353 -680 -352
rect -682 -356 -680 -353
rect -672 -356 -670 -351
rect -664 -353 -660 -351
rect -662 -356 -660 -353
rect -655 -356 -653 -347
rect -614 -351 -612 -343
rect -598 -347 -596 -343
rect -584 -346 -583 -342
rect -579 -346 -578 -342
rect -584 -347 -578 -346
rect -574 -342 -568 -341
rect -574 -346 -573 -342
rect -569 -346 -568 -342
rect -574 -347 -568 -346
rect -544 -342 -542 -339
rect -534 -342 -532 -339
rect -544 -343 -538 -342
rect -544 -347 -543 -343
rect -539 -347 -538 -343
rect -534 -345 -530 -342
rect -605 -348 -596 -347
rect -698 -363 -696 -360
rect -698 -365 -693 -363
rect -764 -373 -762 -368
rect -757 -373 -755 -368
rect -695 -373 -693 -365
rect -682 -369 -680 -365
rect -672 -373 -670 -365
rect -605 -352 -604 -348
rect -600 -352 -596 -348
rect -580 -351 -578 -347
rect -605 -353 -596 -352
rect -598 -356 -596 -353
rect -588 -356 -586 -351
rect -580 -353 -576 -351
rect -578 -356 -576 -353
rect -571 -356 -569 -347
rect -544 -348 -538 -347
rect -544 -356 -542 -348
rect -614 -363 -612 -360
rect -614 -365 -609 -363
rect -662 -373 -660 -368
rect -655 -373 -653 -368
rect -695 -375 -670 -373
rect -611 -373 -609 -365
rect -598 -369 -596 -365
rect -588 -373 -586 -365
rect -532 -359 -530 -345
rect -524 -350 -522 -339
rect -447 -340 -445 -337
rect -437 -340 -435 -337
rect -447 -341 -441 -340
rect -447 -345 -446 -341
rect -442 -345 -441 -341
rect -437 -343 -433 -340
rect -447 -346 -441 -345
rect -525 -351 -519 -350
rect -525 -355 -524 -351
rect -520 -355 -519 -351
rect -447 -354 -445 -346
rect -525 -356 -519 -355
rect -525 -359 -523 -356
rect -544 -366 -542 -362
rect -435 -357 -433 -343
rect -427 -348 -425 -337
rect -372 -339 -370 -330
rect -325 -309 -323 -305
rect -277 -309 -275 -305
rect -345 -318 -343 -314
rect -335 -318 -333 -314
rect -292 -325 -286 -324
rect -292 -329 -291 -325
rect -287 -329 -286 -325
rect -292 -330 -286 -329
rect -361 -339 -359 -336
rect -345 -339 -343 -336
rect -335 -339 -333 -336
rect -325 -339 -323 -336
rect -372 -341 -359 -339
rect -353 -341 -343 -339
rect -339 -340 -333 -339
rect -428 -349 -422 -348
rect -369 -349 -367 -341
rect -353 -345 -351 -341
rect -339 -344 -338 -340
rect -334 -344 -333 -340
rect -339 -345 -333 -344
rect -329 -340 -323 -339
rect -329 -344 -328 -340
rect -324 -344 -323 -340
rect -288 -339 -286 -330
rect -241 -309 -239 -305
rect -261 -318 -259 -314
rect -251 -318 -249 -314
rect -34 -306 -32 -302
rect -110 -314 -104 -313
rect -205 -317 -199 -316
rect -215 -325 -213 -320
rect -205 -321 -204 -317
rect -200 -321 -199 -317
rect -205 -322 -199 -321
rect -120 -322 -118 -317
rect -110 -318 -109 -314
rect -105 -318 -104 -314
rect -110 -319 -104 -318
rect -277 -339 -275 -336
rect -261 -339 -259 -336
rect -251 -339 -249 -336
rect -241 -339 -239 -336
rect -205 -327 -203 -322
rect -195 -327 -193 -322
rect -110 -324 -108 -319
rect -100 -324 -98 -319
rect -49 -322 -43 -321
rect -49 -326 -48 -322
rect -44 -326 -43 -322
rect -49 -327 -43 -326
rect -120 -337 -118 -334
rect -110 -337 -108 -334
rect -288 -341 -275 -339
rect -269 -341 -259 -339
rect -255 -340 -249 -339
rect -329 -345 -323 -344
rect -360 -346 -351 -345
rect -428 -353 -427 -349
rect -423 -353 -422 -349
rect -428 -354 -422 -353
rect -428 -357 -426 -354
rect -447 -364 -445 -360
rect -360 -350 -359 -346
rect -355 -350 -351 -346
rect -335 -349 -333 -345
rect -360 -351 -351 -350
rect -353 -354 -351 -351
rect -343 -354 -341 -349
rect -335 -351 -331 -349
rect -333 -354 -331 -351
rect -326 -354 -324 -345
rect -285 -349 -283 -341
rect -269 -345 -267 -341
rect -255 -344 -254 -340
rect -250 -344 -249 -340
rect -255 -345 -249 -344
rect -245 -340 -239 -339
rect -245 -344 -244 -340
rect -240 -344 -239 -340
rect -245 -345 -239 -344
rect -215 -340 -213 -337
rect -205 -340 -203 -337
rect -215 -341 -209 -340
rect -215 -345 -214 -341
rect -210 -345 -209 -341
rect -205 -343 -201 -340
rect -276 -346 -267 -345
rect -369 -361 -367 -358
rect -369 -363 -364 -361
rect -578 -373 -576 -368
rect -571 -373 -569 -368
rect -611 -375 -586 -373
rect -532 -373 -530 -368
rect -525 -373 -523 -368
rect -435 -371 -433 -366
rect -428 -371 -426 -366
rect -366 -371 -364 -363
rect -353 -367 -351 -363
rect -343 -371 -341 -363
rect -276 -350 -275 -346
rect -271 -350 -267 -346
rect -251 -349 -249 -345
rect -276 -351 -267 -350
rect -269 -354 -267 -351
rect -259 -354 -257 -349
rect -251 -351 -247 -349
rect -249 -354 -247 -351
rect -242 -354 -240 -345
rect -215 -346 -209 -345
rect -215 -354 -213 -346
rect -285 -361 -283 -358
rect -285 -363 -280 -361
rect -333 -371 -331 -366
rect -326 -371 -324 -366
rect -366 -373 -341 -371
rect -282 -371 -280 -363
rect -269 -367 -267 -363
rect -259 -371 -257 -363
rect -203 -357 -201 -343
rect -195 -348 -193 -337
rect -120 -338 -114 -337
rect -120 -342 -119 -338
rect -115 -342 -114 -338
rect -110 -340 -106 -337
rect -120 -343 -114 -342
rect -196 -349 -190 -348
rect -196 -353 -195 -349
rect -191 -353 -190 -349
rect -120 -351 -118 -343
rect -196 -354 -190 -353
rect -196 -357 -194 -354
rect -108 -354 -106 -340
rect -100 -345 -98 -334
rect -45 -336 -43 -327
rect 2 -306 4 -302
rect 50 -306 52 -302
rect -18 -315 -16 -311
rect -8 -315 -6 -311
rect 35 -322 41 -321
rect 35 -326 36 -322
rect 40 -326 41 -322
rect 35 -327 41 -326
rect -34 -336 -32 -333
rect -18 -336 -16 -333
rect -8 -336 -6 -333
rect 2 -336 4 -333
rect -45 -338 -32 -336
rect -26 -338 -16 -336
rect -12 -337 -6 -336
rect -101 -346 -95 -345
rect -42 -346 -40 -338
rect -26 -342 -24 -338
rect -12 -341 -11 -337
rect -7 -341 -6 -337
rect -12 -342 -6 -341
rect -2 -337 4 -336
rect -2 -341 -1 -337
rect 3 -341 4 -337
rect 39 -336 41 -327
rect 86 -306 88 -302
rect 66 -315 68 -311
rect 76 -315 78 -311
rect 122 -314 128 -313
rect 112 -322 114 -317
rect 122 -318 123 -314
rect 127 -318 128 -314
rect 122 -319 128 -318
rect 50 -336 52 -333
rect 66 -336 68 -333
rect 76 -336 78 -333
rect 86 -336 88 -333
rect 122 -324 124 -319
rect 132 -324 134 -319
rect 39 -338 52 -336
rect 58 -338 68 -336
rect 72 -337 78 -336
rect -2 -342 4 -341
rect -33 -343 -24 -342
rect -101 -350 -100 -346
rect -96 -350 -95 -346
rect -101 -351 -95 -350
rect -101 -354 -99 -351
rect -215 -364 -213 -360
rect -120 -361 -118 -357
rect -33 -347 -32 -343
rect -28 -347 -24 -343
rect -8 -346 -6 -342
rect -33 -348 -24 -347
rect -26 -351 -24 -348
rect -16 -351 -14 -346
rect -8 -348 -4 -346
rect -6 -351 -4 -348
rect 1 -351 3 -342
rect 42 -346 44 -338
rect 58 -342 60 -338
rect 72 -341 73 -337
rect 77 -341 78 -337
rect 72 -342 78 -341
rect 82 -337 88 -336
rect 82 -341 83 -337
rect 87 -341 88 -337
rect 82 -342 88 -341
rect 112 -337 114 -334
rect 122 -337 124 -334
rect 112 -338 118 -337
rect 112 -342 113 -338
rect 117 -342 118 -338
rect 122 -340 126 -337
rect 51 -343 60 -342
rect -42 -358 -40 -355
rect -42 -360 -37 -358
rect -249 -371 -247 -366
rect -242 -371 -240 -366
rect -282 -373 -257 -371
rect -203 -371 -201 -366
rect -196 -371 -194 -366
rect -108 -368 -106 -363
rect -101 -368 -99 -363
rect -39 -368 -37 -360
rect -26 -364 -24 -360
rect -16 -368 -14 -360
rect 51 -347 52 -343
rect 56 -347 60 -343
rect 76 -346 78 -342
rect 51 -348 60 -347
rect 58 -351 60 -348
rect 68 -351 70 -346
rect 76 -348 80 -346
rect 78 -351 80 -348
rect 85 -351 87 -342
rect 112 -343 118 -342
rect 112 -351 114 -343
rect 42 -358 44 -355
rect 42 -360 47 -358
rect -6 -368 -4 -363
rect 1 -368 3 -363
rect -39 -370 -14 -368
rect 45 -368 47 -360
rect 58 -364 60 -360
rect 68 -368 70 -360
rect 124 -354 126 -340
rect 132 -345 134 -334
rect 131 -346 137 -345
rect 131 -350 132 -346
rect 136 -350 137 -346
rect 131 -351 137 -350
rect 131 -354 133 -351
rect 112 -361 114 -357
rect 78 -368 80 -363
rect 85 -368 87 -363
rect 45 -370 70 -368
rect 124 -368 126 -363
rect 131 -368 133 -363
rect -683 -390 -681 -386
rect -673 -390 -671 -386
rect -663 -390 -661 -386
rect -354 -388 -352 -384
rect -344 -388 -342 -384
rect -334 -388 -332 -384
rect -27 -385 -25 -381
rect -17 -385 -15 -381
rect -7 -385 -5 -381
rect -683 -404 -681 -396
rect -687 -405 -681 -404
rect -673 -405 -671 -396
rect -663 -405 -661 -396
rect -354 -402 -352 -394
rect -687 -409 -686 -405
rect -682 -409 -681 -405
rect -667 -406 -661 -405
rect -687 -410 -681 -409
rect -683 -423 -681 -410
rect -673 -412 -671 -409
rect -667 -410 -666 -406
rect -662 -410 -661 -406
rect -358 -403 -352 -402
rect -344 -403 -342 -394
rect -334 -403 -332 -394
rect -27 -399 -25 -391
rect -358 -407 -357 -403
rect -353 -407 -352 -403
rect -338 -404 -332 -403
rect -358 -408 -352 -407
rect -667 -411 -661 -410
rect -677 -413 -671 -412
rect -677 -417 -676 -413
rect -672 -417 -671 -413
rect -677 -418 -671 -417
rect -676 -423 -674 -418
rect -663 -420 -661 -411
rect -354 -421 -352 -408
rect -344 -410 -342 -407
rect -338 -408 -337 -404
rect -333 -408 -332 -404
rect -31 -400 -25 -399
rect -17 -400 -15 -391
rect -7 -400 -5 -391
rect -31 -404 -30 -400
rect -26 -404 -25 -400
rect -11 -401 -5 -400
rect -31 -405 -25 -404
rect -338 -409 -332 -408
rect -348 -411 -342 -410
rect -348 -415 -347 -411
rect -343 -415 -342 -411
rect -348 -416 -342 -415
rect -347 -421 -345 -416
rect -334 -418 -332 -409
rect -27 -418 -25 -405
rect -17 -407 -15 -404
rect -11 -405 -10 -401
rect -6 -405 -5 -401
rect -11 -406 -5 -405
rect -21 -408 -15 -407
rect -21 -412 -20 -408
rect -16 -412 -15 -408
rect -21 -413 -15 -412
rect -20 -418 -18 -413
rect -7 -415 -5 -406
rect -663 -436 -661 -432
rect -334 -434 -332 -430
rect -7 -431 -5 -427
rect -683 -445 -681 -441
rect -676 -445 -674 -441
rect -354 -443 -352 -439
rect -347 -443 -345 -439
rect -27 -440 -25 -436
rect -20 -440 -18 -436
rect -482 -468 -480 -464
rect -472 -466 -470 -461
rect -462 -466 -460 -461
rect -389 -468 -387 -464
rect -379 -466 -377 -461
rect -369 -466 -367 -461
rect -482 -490 -480 -486
rect -472 -490 -470 -479
rect -462 -482 -460 -479
rect -462 -483 -456 -482
rect -462 -487 -461 -483
rect -457 -487 -456 -483
rect -302 -468 -300 -464
rect -292 -466 -290 -461
rect -282 -466 -280 -461
rect -462 -488 -456 -487
rect -482 -491 -476 -490
rect -482 -495 -481 -491
rect -477 -495 -476 -491
rect -482 -496 -476 -495
rect -472 -491 -466 -490
rect -472 -495 -471 -491
rect -467 -495 -466 -491
rect -472 -496 -466 -495
rect -482 -501 -480 -496
rect -469 -501 -467 -496
rect -462 -501 -460 -488
rect -389 -490 -387 -486
rect -379 -490 -377 -479
rect -369 -482 -367 -479
rect -369 -483 -363 -482
rect -369 -487 -368 -483
rect -364 -487 -363 -483
rect -369 -488 -363 -487
rect -389 -491 -383 -490
rect -389 -495 -388 -491
rect -384 -495 -383 -491
rect -389 -496 -383 -495
rect -379 -491 -373 -490
rect -379 -495 -378 -491
rect -374 -495 -373 -491
rect -379 -496 -373 -495
rect -389 -501 -387 -496
rect -376 -501 -374 -496
rect -369 -501 -367 -488
rect -302 -490 -300 -486
rect -292 -490 -290 -479
rect -282 -482 -280 -479
rect -282 -483 -276 -482
rect -282 -487 -281 -483
rect -277 -487 -276 -483
rect -282 -488 -276 -487
rect -302 -491 -296 -490
rect -302 -495 -301 -491
rect -297 -495 -296 -491
rect -302 -496 -296 -495
rect -292 -491 -286 -490
rect -292 -495 -291 -491
rect -287 -495 -286 -491
rect -292 -496 -286 -495
rect -302 -501 -300 -496
rect -289 -501 -287 -496
rect -282 -501 -280 -488
rect -482 -514 -480 -510
rect -469 -517 -467 -512
rect -462 -517 -460 -512
rect -389 -514 -387 -510
rect -376 -517 -374 -512
rect -369 -517 -367 -512
rect -302 -514 -300 -510
rect -289 -517 -287 -512
rect -282 -517 -280 -512
<< ndiffusion >>
rect -89 -71 -78 -68
rect -76 -71 -59 -68
rect 23 -67 33 -66
rect -17 -72 -6 -69
rect -4 -72 13 -69
rect 23 -71 25 -67
rect 29 -71 33 -67
rect 23 -72 33 -71
rect 35 -72 54 -66
rect 56 -67 64 -66
rect 56 -71 59 -67
rect 63 -71 64 -67
rect 56 -72 64 -71
rect 77 -67 87 -66
rect 77 -71 79 -67
rect 83 -71 87 -67
rect 77 -72 87 -71
rect 89 -72 108 -66
rect 110 -67 118 -66
rect 110 -71 113 -67
rect 117 -71 118 -67
rect 110 -72 118 -71
rect 133 -67 143 -66
rect 133 -71 135 -67
rect 139 -71 143 -67
rect 133 -72 143 -71
rect 145 -72 164 -66
rect 166 -67 174 -66
rect 166 -71 169 -67
rect 173 -71 174 -67
rect 166 -72 174 -71
rect 187 -67 197 -66
rect 187 -71 189 -67
rect 193 -71 197 -67
rect 187 -72 197 -71
rect 199 -72 218 -66
rect 220 -67 228 -66
rect 220 -71 223 -67
rect 227 -71 228 -67
rect 220 -72 228 -71
rect -686 -84 -679 -83
rect -686 -88 -684 -84
rect -680 -88 -679 -84
rect -686 -93 -679 -88
rect -599 -84 -592 -83
rect -599 -88 -597 -84
rect -593 -88 -592 -84
rect -704 -94 -697 -93
rect -704 -98 -703 -94
rect -699 -98 -697 -94
rect -704 -99 -697 -98
rect -702 -104 -697 -99
rect -695 -104 -690 -93
rect -688 -95 -679 -93
rect -599 -93 -592 -88
rect -506 -84 -499 -83
rect -506 -88 -504 -84
rect -500 -88 -499 -84
rect -617 -94 -610 -93
rect -688 -104 -677 -95
rect -675 -96 -668 -95
rect -675 -100 -673 -96
rect -669 -100 -668 -96
rect -617 -98 -616 -94
rect -612 -98 -610 -94
rect -617 -99 -610 -98
rect -675 -101 -668 -100
rect -675 -104 -670 -101
rect -615 -104 -610 -99
rect -608 -104 -603 -93
rect -601 -95 -592 -93
rect -506 -93 -499 -88
rect -273 -82 -266 -81
rect -273 -86 -272 -82
rect -268 -86 -266 -82
rect -524 -94 -517 -93
rect -601 -104 -590 -95
rect -588 -96 -581 -95
rect -588 -100 -586 -96
rect -582 -100 -581 -96
rect -524 -98 -523 -94
rect -519 -98 -517 -94
rect -524 -99 -517 -98
rect -588 -101 -581 -100
rect -588 -104 -583 -101
rect -522 -104 -517 -99
rect -515 -104 -510 -93
rect -508 -95 -499 -93
rect -273 -91 -266 -86
rect -180 -82 -173 -81
rect -180 -86 -179 -82
rect -175 -86 -173 -82
rect -273 -93 -264 -91
rect -284 -94 -277 -93
rect -508 -104 -497 -95
rect -495 -96 -488 -95
rect -495 -100 -493 -96
rect -489 -100 -488 -96
rect -284 -98 -283 -94
rect -279 -98 -277 -94
rect -284 -99 -277 -98
rect -495 -101 -488 -100
rect -495 -104 -490 -101
rect -282 -102 -277 -99
rect -275 -102 -264 -93
rect -262 -102 -257 -91
rect -255 -92 -248 -91
rect -255 -96 -253 -92
rect -249 -96 -248 -92
rect -180 -91 -173 -86
rect -93 -82 -86 -81
rect -93 -86 -92 -82
rect -88 -86 -86 -82
rect -180 -93 -171 -91
rect -255 -97 -248 -96
rect -191 -94 -184 -93
rect -255 -102 -250 -97
rect -191 -98 -190 -94
rect -186 -98 -184 -94
rect -191 -99 -184 -98
rect -189 -102 -184 -99
rect -182 -102 -171 -93
rect -169 -102 -164 -91
rect -162 -92 -155 -91
rect -162 -96 -160 -92
rect -156 -96 -155 -92
rect -93 -91 -86 -86
rect -93 -93 -84 -91
rect -162 -97 -155 -96
rect -104 -94 -97 -93
rect -162 -102 -157 -97
rect -104 -98 -103 -94
rect -99 -98 -97 -94
rect -104 -99 -97 -98
rect -102 -102 -97 -99
rect -95 -102 -84 -93
rect -82 -102 -77 -91
rect -75 -92 -68 -91
rect -75 -96 -73 -92
rect -69 -96 -68 -92
rect -13 -94 -2 -91
rect 0 -94 17 -91
rect -75 -97 -68 -96
rect -75 -102 -70 -97
rect 27 -92 37 -91
rect 27 -96 29 -92
rect 33 -96 37 -92
rect 27 -97 37 -96
rect 39 -97 58 -91
rect 60 -92 68 -91
rect 60 -96 63 -92
rect 67 -96 68 -92
rect 60 -97 68 -96
rect 81 -92 91 -91
rect 81 -96 83 -92
rect 87 -96 91 -92
rect 81 -97 91 -96
rect 93 -97 112 -91
rect 114 -92 122 -91
rect 114 -96 117 -92
rect 121 -96 122 -92
rect 114 -97 122 -96
rect 137 -92 147 -91
rect 137 -96 139 -92
rect 143 -96 147 -92
rect 137 -97 147 -96
rect 149 -97 168 -91
rect 170 -92 178 -91
rect 170 -96 173 -92
rect 177 -96 178 -92
rect 170 -97 178 -96
rect 191 -92 201 -91
rect 191 -96 193 -92
rect 197 -96 201 -92
rect 191 -97 201 -96
rect 203 -97 222 -91
rect 224 -92 232 -91
rect 224 -96 227 -92
rect 231 -96 232 -92
rect 224 -97 232 -96
rect -782 -211 -775 -210
rect -782 -215 -781 -211
rect -777 -215 -775 -211
rect -782 -216 -775 -215
rect -773 -213 -765 -210
rect -704 -206 -697 -205
rect -704 -210 -703 -206
rect -699 -210 -697 -206
rect -704 -211 -697 -210
rect -773 -216 -763 -213
rect -771 -222 -763 -216
rect -761 -222 -756 -213
rect -754 -214 -747 -213
rect -702 -214 -697 -211
rect -695 -210 -690 -205
rect -620 -206 -613 -205
rect -620 -210 -619 -206
rect -615 -210 -613 -206
rect -695 -214 -681 -210
rect -754 -218 -752 -214
rect -748 -218 -747 -214
rect -754 -219 -747 -218
rect -690 -218 -689 -214
rect -685 -218 -681 -214
rect -690 -219 -681 -218
rect -679 -211 -671 -210
rect -679 -215 -677 -211
rect -673 -215 -671 -211
rect -679 -219 -671 -215
rect -669 -213 -661 -210
rect -669 -217 -667 -213
rect -663 -217 -661 -213
rect -669 -219 -661 -217
rect -754 -222 -749 -219
rect -771 -223 -765 -222
rect -771 -227 -770 -223
rect -766 -227 -765 -223
rect -771 -228 -765 -227
rect -666 -222 -661 -219
rect -659 -222 -654 -210
rect -652 -222 -644 -210
rect -620 -211 -613 -210
rect -618 -214 -613 -211
rect -611 -210 -606 -205
rect -611 -214 -597 -210
rect -606 -218 -605 -214
rect -601 -218 -597 -214
rect -606 -219 -597 -218
rect -595 -211 -587 -210
rect -595 -215 -593 -211
rect -589 -215 -587 -211
rect -595 -219 -587 -215
rect -585 -213 -577 -210
rect -585 -217 -583 -213
rect -579 -217 -577 -213
rect -585 -219 -577 -217
rect -650 -223 -644 -222
rect -650 -227 -649 -223
rect -645 -227 -644 -223
rect -650 -228 -644 -227
rect -582 -222 -577 -219
rect -575 -222 -570 -210
rect -568 -222 -560 -210
rect -550 -211 -543 -210
rect -550 -215 -549 -211
rect -545 -215 -543 -211
rect -550 -216 -543 -215
rect -541 -213 -533 -210
rect -453 -209 -446 -208
rect -453 -213 -452 -209
rect -448 -213 -446 -209
rect -541 -216 -531 -213
rect -539 -222 -531 -216
rect -529 -222 -524 -213
rect -522 -214 -515 -213
rect -453 -214 -446 -213
rect -444 -211 -436 -208
rect -375 -204 -368 -203
rect -375 -208 -374 -204
rect -370 -208 -368 -204
rect -375 -209 -368 -208
rect -444 -214 -434 -211
rect -522 -218 -520 -214
rect -516 -218 -515 -214
rect -522 -219 -515 -218
rect -522 -222 -517 -219
rect -442 -220 -434 -214
rect -432 -220 -427 -211
rect -425 -212 -418 -211
rect -373 -212 -368 -209
rect -366 -208 -361 -203
rect -291 -204 -284 -203
rect -291 -208 -290 -204
rect -286 -208 -284 -204
rect -366 -212 -352 -208
rect -425 -216 -423 -212
rect -419 -216 -418 -212
rect -425 -217 -418 -216
rect -361 -216 -360 -212
rect -356 -216 -352 -212
rect -361 -217 -352 -216
rect -350 -209 -342 -208
rect -350 -213 -348 -209
rect -344 -213 -342 -209
rect -350 -217 -342 -213
rect -340 -211 -332 -208
rect -340 -215 -338 -211
rect -334 -215 -332 -211
rect -340 -217 -332 -215
rect -425 -220 -420 -217
rect -566 -223 -560 -222
rect -566 -227 -565 -223
rect -561 -227 -560 -223
rect -566 -228 -560 -227
rect -539 -223 -533 -222
rect -539 -227 -538 -223
rect -534 -227 -533 -223
rect -442 -221 -436 -220
rect -442 -225 -441 -221
rect -437 -225 -436 -221
rect -442 -226 -436 -225
rect -337 -220 -332 -217
rect -330 -220 -325 -208
rect -323 -220 -315 -208
rect -291 -209 -284 -208
rect -289 -212 -284 -209
rect -282 -208 -277 -203
rect -282 -212 -268 -208
rect -277 -216 -276 -212
rect -272 -216 -268 -212
rect -277 -217 -268 -216
rect -266 -209 -258 -208
rect -266 -213 -264 -209
rect -260 -213 -258 -209
rect -266 -217 -258 -213
rect -256 -211 -248 -208
rect -256 -215 -254 -211
rect -250 -215 -248 -211
rect -256 -217 -248 -215
rect -321 -221 -315 -220
rect -321 -225 -320 -221
rect -316 -225 -315 -221
rect -321 -226 -315 -225
rect -253 -220 -248 -217
rect -246 -220 -241 -208
rect -239 -220 -231 -208
rect -221 -209 -214 -208
rect -221 -213 -220 -209
rect -216 -213 -214 -209
rect -221 -214 -214 -213
rect -212 -211 -204 -208
rect -126 -206 -119 -205
rect -126 -210 -125 -206
rect -121 -210 -119 -206
rect -126 -211 -119 -210
rect -117 -208 -109 -205
rect -48 -201 -41 -200
rect -48 -205 -47 -201
rect -43 -205 -41 -201
rect -48 -206 -41 -205
rect -117 -211 -107 -208
rect -212 -214 -202 -211
rect -210 -220 -202 -214
rect -200 -220 -195 -211
rect -193 -212 -186 -211
rect -193 -216 -191 -212
rect -187 -216 -186 -212
rect -193 -217 -186 -216
rect -115 -217 -107 -211
rect -105 -217 -100 -208
rect -98 -209 -91 -208
rect -46 -209 -41 -206
rect -39 -205 -34 -200
rect 36 -201 43 -200
rect 36 -205 37 -201
rect 41 -205 43 -201
rect -39 -209 -25 -205
rect -98 -213 -96 -209
rect -92 -213 -91 -209
rect -98 -214 -91 -213
rect -34 -213 -33 -209
rect -29 -213 -25 -209
rect -34 -214 -25 -213
rect -23 -206 -15 -205
rect -23 -210 -21 -206
rect -17 -210 -15 -206
rect -23 -214 -15 -210
rect -13 -208 -5 -205
rect -13 -212 -11 -208
rect -7 -212 -5 -208
rect -13 -214 -5 -212
rect -98 -217 -93 -214
rect -193 -220 -188 -217
rect -237 -221 -231 -220
rect -237 -225 -236 -221
rect -232 -225 -231 -221
rect -237 -226 -231 -225
rect -210 -221 -204 -220
rect -210 -225 -209 -221
rect -205 -225 -204 -221
rect -115 -218 -109 -217
rect -115 -222 -114 -218
rect -110 -222 -109 -218
rect -115 -223 -109 -222
rect -10 -217 -5 -214
rect -3 -217 2 -205
rect 4 -217 12 -205
rect 36 -206 43 -205
rect 38 -209 43 -206
rect 45 -205 50 -200
rect 45 -209 59 -205
rect 50 -213 51 -209
rect 55 -213 59 -209
rect 50 -214 59 -213
rect 61 -206 69 -205
rect 61 -210 63 -206
rect 67 -210 69 -206
rect 61 -214 69 -210
rect 71 -208 79 -205
rect 71 -212 73 -208
rect 77 -212 79 -208
rect 71 -214 79 -212
rect 6 -218 12 -217
rect 6 -222 7 -218
rect 11 -222 12 -218
rect 6 -223 12 -222
rect 74 -217 79 -214
rect 81 -217 86 -205
rect 88 -217 96 -205
rect 106 -206 113 -205
rect 106 -210 107 -206
rect 111 -210 113 -206
rect 106 -211 113 -210
rect 115 -208 123 -205
rect 115 -211 125 -208
rect 117 -217 125 -211
rect 127 -217 132 -208
rect 134 -209 141 -208
rect 134 -213 136 -209
rect 140 -213 141 -209
rect 134 -214 141 -213
rect 134 -217 139 -214
rect 90 -218 96 -217
rect 90 -222 91 -218
rect 95 -222 96 -218
rect 90 -223 96 -222
rect 117 -218 123 -217
rect 117 -222 118 -218
rect 122 -222 123 -218
rect 117 -223 123 -222
rect -210 -226 -204 -225
rect -539 -228 -533 -227
rect -33 -240 -26 -239
rect -360 -243 -353 -242
rect -689 -245 -682 -244
rect -689 -249 -688 -245
rect -684 -249 -682 -245
rect -689 -250 -682 -249
rect -680 -245 -672 -244
rect -680 -249 -678 -245
rect -674 -249 -672 -245
rect -680 -250 -672 -249
rect -670 -245 -662 -244
rect -670 -249 -668 -245
rect -664 -249 -662 -245
rect -670 -250 -662 -249
rect -660 -245 -653 -244
rect -660 -249 -658 -245
rect -654 -249 -653 -245
rect -360 -247 -359 -243
rect -355 -247 -353 -243
rect -360 -248 -353 -247
rect -351 -243 -343 -242
rect -351 -247 -349 -243
rect -345 -247 -343 -243
rect -351 -248 -343 -247
rect -341 -243 -333 -242
rect -341 -247 -339 -243
rect -335 -247 -333 -243
rect -341 -248 -333 -247
rect -331 -243 -324 -242
rect -331 -247 -329 -243
rect -325 -247 -324 -243
rect -33 -244 -32 -240
rect -28 -244 -26 -240
rect -33 -245 -26 -244
rect -24 -240 -16 -239
rect -24 -244 -22 -240
rect -18 -244 -16 -240
rect -24 -245 -16 -244
rect -14 -240 -6 -239
rect -14 -244 -12 -240
rect -8 -244 -6 -240
rect -14 -245 -6 -244
rect -4 -240 3 -239
rect -4 -244 -2 -240
rect 2 -244 3 -240
rect -4 -245 3 -244
rect -331 -248 -324 -247
rect -660 -250 -653 -249
rect -783 -357 -776 -356
rect -783 -361 -782 -357
rect -778 -361 -776 -357
rect -783 -362 -776 -361
rect -774 -359 -766 -356
rect -705 -352 -698 -351
rect -705 -356 -704 -352
rect -700 -356 -698 -352
rect -705 -357 -698 -356
rect -774 -362 -764 -359
rect -772 -368 -764 -362
rect -762 -368 -757 -359
rect -755 -360 -748 -359
rect -703 -360 -698 -357
rect -696 -356 -691 -351
rect -621 -352 -614 -351
rect -621 -356 -620 -352
rect -616 -356 -614 -352
rect -696 -360 -682 -356
rect -755 -364 -753 -360
rect -749 -364 -748 -360
rect -755 -365 -748 -364
rect -691 -364 -690 -360
rect -686 -364 -682 -360
rect -691 -365 -682 -364
rect -680 -357 -672 -356
rect -680 -361 -678 -357
rect -674 -361 -672 -357
rect -680 -365 -672 -361
rect -670 -359 -662 -356
rect -670 -363 -668 -359
rect -664 -363 -662 -359
rect -670 -365 -662 -363
rect -755 -368 -750 -365
rect -772 -369 -766 -368
rect -772 -373 -771 -369
rect -767 -373 -766 -369
rect -772 -374 -766 -373
rect -667 -368 -662 -365
rect -660 -368 -655 -356
rect -653 -368 -645 -356
rect -621 -357 -614 -356
rect -619 -360 -614 -357
rect -612 -356 -607 -351
rect -612 -360 -598 -356
rect -607 -364 -606 -360
rect -602 -364 -598 -360
rect -607 -365 -598 -364
rect -596 -357 -588 -356
rect -596 -361 -594 -357
rect -590 -361 -588 -357
rect -596 -365 -588 -361
rect -586 -359 -578 -356
rect -586 -363 -584 -359
rect -580 -363 -578 -359
rect -586 -365 -578 -363
rect -651 -369 -645 -368
rect -651 -373 -650 -369
rect -646 -373 -645 -369
rect -651 -374 -645 -373
rect -583 -368 -578 -365
rect -576 -368 -571 -356
rect -569 -368 -561 -356
rect -551 -357 -544 -356
rect -551 -361 -550 -357
rect -546 -361 -544 -357
rect -551 -362 -544 -361
rect -542 -359 -534 -356
rect -454 -355 -447 -354
rect -454 -359 -453 -355
rect -449 -359 -447 -355
rect -542 -362 -532 -359
rect -540 -368 -532 -362
rect -530 -368 -525 -359
rect -523 -360 -516 -359
rect -454 -360 -447 -359
rect -445 -357 -437 -354
rect -376 -350 -369 -349
rect -376 -354 -375 -350
rect -371 -354 -369 -350
rect -376 -355 -369 -354
rect -445 -360 -435 -357
rect -523 -364 -521 -360
rect -517 -364 -516 -360
rect -523 -365 -516 -364
rect -523 -368 -518 -365
rect -443 -366 -435 -360
rect -433 -366 -428 -357
rect -426 -358 -419 -357
rect -374 -358 -369 -355
rect -367 -354 -362 -349
rect -292 -350 -285 -349
rect -292 -354 -291 -350
rect -287 -354 -285 -350
rect -367 -358 -353 -354
rect -426 -362 -424 -358
rect -420 -362 -419 -358
rect -426 -363 -419 -362
rect -362 -362 -361 -358
rect -357 -362 -353 -358
rect -362 -363 -353 -362
rect -351 -355 -343 -354
rect -351 -359 -349 -355
rect -345 -359 -343 -355
rect -351 -363 -343 -359
rect -341 -357 -333 -354
rect -341 -361 -339 -357
rect -335 -361 -333 -357
rect -341 -363 -333 -361
rect -426 -366 -421 -363
rect -567 -369 -561 -368
rect -567 -373 -566 -369
rect -562 -373 -561 -369
rect -567 -374 -561 -373
rect -540 -369 -534 -368
rect -540 -373 -539 -369
rect -535 -373 -534 -369
rect -443 -367 -437 -366
rect -443 -371 -442 -367
rect -438 -371 -437 -367
rect -443 -372 -437 -371
rect -338 -366 -333 -363
rect -331 -366 -326 -354
rect -324 -366 -316 -354
rect -292 -355 -285 -354
rect -290 -358 -285 -355
rect -283 -354 -278 -349
rect -283 -358 -269 -354
rect -278 -362 -277 -358
rect -273 -362 -269 -358
rect -278 -363 -269 -362
rect -267 -355 -259 -354
rect -267 -359 -265 -355
rect -261 -359 -259 -355
rect -267 -363 -259 -359
rect -257 -357 -249 -354
rect -257 -361 -255 -357
rect -251 -361 -249 -357
rect -257 -363 -249 -361
rect -322 -367 -316 -366
rect -322 -371 -321 -367
rect -317 -371 -316 -367
rect -322 -372 -316 -371
rect -254 -366 -249 -363
rect -247 -366 -242 -354
rect -240 -366 -232 -354
rect -222 -355 -215 -354
rect -222 -359 -221 -355
rect -217 -359 -215 -355
rect -222 -360 -215 -359
rect -213 -357 -205 -354
rect -127 -352 -120 -351
rect -127 -356 -126 -352
rect -122 -356 -120 -352
rect -127 -357 -120 -356
rect -118 -354 -110 -351
rect -49 -347 -42 -346
rect -49 -351 -48 -347
rect -44 -351 -42 -347
rect -49 -352 -42 -351
rect -118 -357 -108 -354
rect -213 -360 -203 -357
rect -211 -366 -203 -360
rect -201 -366 -196 -357
rect -194 -358 -187 -357
rect -194 -362 -192 -358
rect -188 -362 -187 -358
rect -194 -363 -187 -362
rect -116 -363 -108 -357
rect -106 -363 -101 -354
rect -99 -355 -92 -354
rect -47 -355 -42 -352
rect -40 -351 -35 -346
rect 35 -347 42 -346
rect 35 -351 36 -347
rect 40 -351 42 -347
rect -40 -355 -26 -351
rect -99 -359 -97 -355
rect -93 -359 -92 -355
rect -99 -360 -92 -359
rect -35 -359 -34 -355
rect -30 -359 -26 -355
rect -35 -360 -26 -359
rect -24 -352 -16 -351
rect -24 -356 -22 -352
rect -18 -356 -16 -352
rect -24 -360 -16 -356
rect -14 -354 -6 -351
rect -14 -358 -12 -354
rect -8 -358 -6 -354
rect -14 -360 -6 -358
rect -99 -363 -94 -360
rect -194 -366 -189 -363
rect -238 -367 -232 -366
rect -238 -371 -237 -367
rect -233 -371 -232 -367
rect -238 -372 -232 -371
rect -211 -367 -205 -366
rect -211 -371 -210 -367
rect -206 -371 -205 -367
rect -116 -364 -110 -363
rect -116 -368 -115 -364
rect -111 -368 -110 -364
rect -116 -369 -110 -368
rect -11 -363 -6 -360
rect -4 -363 1 -351
rect 3 -363 11 -351
rect 35 -352 42 -351
rect 37 -355 42 -352
rect 44 -351 49 -346
rect 44 -355 58 -351
rect 49 -359 50 -355
rect 54 -359 58 -355
rect 49 -360 58 -359
rect 60 -352 68 -351
rect 60 -356 62 -352
rect 66 -356 68 -352
rect 60 -360 68 -356
rect 70 -354 78 -351
rect 70 -358 72 -354
rect 76 -358 78 -354
rect 70 -360 78 -358
rect 5 -364 11 -363
rect 5 -368 6 -364
rect 10 -368 11 -364
rect 5 -369 11 -368
rect 73 -363 78 -360
rect 80 -363 85 -351
rect 87 -363 95 -351
rect 105 -352 112 -351
rect 105 -356 106 -352
rect 110 -356 112 -352
rect 105 -357 112 -356
rect 114 -354 122 -351
rect 114 -357 124 -354
rect 116 -363 124 -357
rect 126 -363 131 -354
rect 133 -355 140 -354
rect 133 -359 135 -355
rect 139 -359 140 -355
rect 133 -360 140 -359
rect 133 -363 138 -360
rect 89 -364 95 -363
rect 89 -368 90 -364
rect 94 -368 95 -364
rect 89 -369 95 -368
rect 116 -364 122 -363
rect 116 -368 117 -364
rect 121 -368 122 -364
rect 116 -369 122 -368
rect -211 -372 -205 -371
rect -540 -374 -534 -373
rect -34 -386 -27 -385
rect -361 -389 -354 -388
rect -690 -391 -683 -390
rect -690 -395 -689 -391
rect -685 -395 -683 -391
rect -690 -396 -683 -395
rect -681 -391 -673 -390
rect -681 -395 -679 -391
rect -675 -395 -673 -391
rect -681 -396 -673 -395
rect -671 -391 -663 -390
rect -671 -395 -669 -391
rect -665 -395 -663 -391
rect -671 -396 -663 -395
rect -661 -391 -654 -390
rect -661 -395 -659 -391
rect -655 -395 -654 -391
rect -361 -393 -360 -389
rect -356 -393 -354 -389
rect -361 -394 -354 -393
rect -352 -389 -344 -388
rect -352 -393 -350 -389
rect -346 -393 -344 -389
rect -352 -394 -344 -393
rect -342 -389 -334 -388
rect -342 -393 -340 -389
rect -336 -393 -334 -389
rect -342 -394 -334 -393
rect -332 -389 -325 -388
rect -332 -393 -330 -389
rect -326 -393 -325 -389
rect -34 -390 -33 -386
rect -29 -390 -27 -386
rect -34 -391 -27 -390
rect -25 -386 -17 -385
rect -25 -390 -23 -386
rect -19 -390 -17 -386
rect -25 -391 -17 -390
rect -15 -386 -7 -385
rect -15 -390 -13 -386
rect -9 -390 -7 -386
rect -15 -391 -7 -390
rect -5 -386 2 -385
rect -5 -390 -3 -386
rect 1 -390 2 -386
rect -5 -391 2 -390
rect -332 -394 -325 -393
rect -661 -396 -654 -395
rect -487 -504 -482 -501
rect -489 -505 -482 -504
rect -489 -509 -488 -505
rect -484 -509 -482 -505
rect -489 -510 -482 -509
rect -480 -510 -469 -501
rect -478 -512 -469 -510
rect -467 -512 -462 -501
rect -460 -506 -455 -501
rect -394 -504 -389 -501
rect -396 -505 -389 -504
rect -460 -507 -453 -506
rect -460 -511 -458 -507
rect -454 -511 -453 -507
rect -396 -509 -395 -505
rect -391 -509 -389 -505
rect -396 -510 -389 -509
rect -387 -510 -376 -501
rect -460 -512 -453 -511
rect -478 -517 -471 -512
rect -385 -512 -376 -510
rect -374 -512 -369 -501
rect -367 -506 -362 -501
rect -307 -504 -302 -501
rect -309 -505 -302 -504
rect -367 -507 -360 -506
rect -367 -511 -365 -507
rect -361 -511 -360 -507
rect -309 -509 -308 -505
rect -304 -509 -302 -505
rect -309 -510 -302 -509
rect -300 -510 -289 -501
rect -367 -512 -360 -511
rect -478 -521 -477 -517
rect -473 -521 -471 -517
rect -478 -522 -471 -521
rect -385 -517 -378 -512
rect -298 -512 -289 -510
rect -287 -512 -282 -501
rect -280 -506 -275 -501
rect -280 -507 -273 -506
rect -280 -511 -278 -507
rect -274 -511 -273 -507
rect -280 -512 -273 -511
rect -385 -521 -384 -517
rect -380 -521 -378 -517
rect -385 -522 -378 -521
rect -298 -517 -291 -512
rect -298 -521 -297 -517
rect -293 -521 -291 -517
rect -298 -522 -291 -521
<< pdiffusion >>
rect -109 -30 -78 -29
rect -109 -34 -104 -30
rect -100 -34 -78 -30
rect -109 -35 -78 -34
rect -76 -34 -60 -29
rect -54 -34 -41 -29
rect -76 -35 -41 -34
rect -21 -30 -6 -29
rect -17 -34 -6 -30
rect -21 -35 -6 -34
rect -4 -30 16 -29
rect -4 -34 12 -30
rect -4 -35 16 -34
rect 23 -30 33 -29
rect 23 -34 25 -30
rect 29 -34 33 -30
rect 23 -35 33 -34
rect 35 -30 54 -29
rect 35 -34 42 -30
rect 46 -34 54 -30
rect 35 -35 54 -34
rect 56 -30 64 -29
rect 56 -34 59 -30
rect 63 -34 64 -30
rect 56 -35 64 -34
rect 77 -30 87 -29
rect 77 -34 79 -30
rect 83 -34 87 -30
rect 77 -35 87 -34
rect 89 -30 108 -29
rect 89 -34 96 -30
rect 100 -34 108 -30
rect 89 -35 108 -34
rect 110 -30 118 -29
rect 110 -34 113 -30
rect 117 -34 118 -30
rect 110 -35 118 -34
rect 133 -30 143 -29
rect 133 -34 135 -30
rect 139 -34 143 -30
rect 133 -35 143 -34
rect 145 -30 164 -29
rect 145 -34 152 -30
rect 156 -34 164 -30
rect 145 -35 164 -34
rect 166 -30 174 -29
rect 166 -34 169 -30
rect 173 -34 174 -30
rect 166 -35 174 -34
rect 187 -30 197 -29
rect 187 -34 189 -30
rect 193 -34 197 -30
rect 187 -35 197 -34
rect 199 -30 218 -29
rect 199 -34 206 -30
rect 210 -34 218 -30
rect 199 -35 218 -34
rect 220 -30 228 -29
rect 220 -34 223 -30
rect 227 -34 228 -30
rect 220 -35 228 -34
rect -683 -126 -677 -119
rect -704 -134 -697 -126
rect -704 -138 -703 -134
rect -699 -138 -697 -134
rect -704 -139 -697 -138
rect -695 -127 -687 -126
rect -695 -131 -693 -127
rect -689 -131 -687 -127
rect -695 -134 -687 -131
rect -695 -138 -693 -134
rect -689 -138 -687 -134
rect -695 -139 -687 -138
rect -685 -132 -677 -126
rect -685 -136 -683 -132
rect -679 -136 -677 -132
rect -685 -137 -677 -136
rect -675 -120 -668 -119
rect -675 -124 -673 -120
rect -669 -124 -668 -120
rect -675 -127 -668 -124
rect -596 -126 -590 -119
rect -675 -131 -673 -127
rect -669 -131 -668 -127
rect -675 -132 -668 -131
rect -675 -137 -670 -132
rect -617 -134 -610 -126
rect -685 -139 -679 -137
rect -617 -138 -616 -134
rect -612 -138 -610 -134
rect -617 -139 -610 -138
rect -608 -127 -600 -126
rect -608 -131 -606 -127
rect -602 -131 -600 -127
rect -608 -134 -600 -131
rect -608 -138 -606 -134
rect -602 -138 -600 -134
rect -608 -139 -600 -138
rect -598 -132 -590 -126
rect -598 -136 -596 -132
rect -592 -136 -590 -132
rect -598 -137 -590 -136
rect -588 -120 -581 -119
rect -588 -124 -586 -120
rect -582 -124 -581 -120
rect -588 -127 -581 -124
rect -284 -118 -277 -117
rect -503 -126 -497 -119
rect -588 -131 -586 -127
rect -582 -131 -581 -127
rect -588 -132 -581 -131
rect -588 -137 -583 -132
rect -524 -134 -517 -126
rect -598 -139 -592 -137
rect -524 -138 -523 -134
rect -519 -138 -517 -134
rect -524 -139 -517 -138
rect -515 -127 -507 -126
rect -515 -131 -513 -127
rect -509 -131 -507 -127
rect -515 -134 -507 -131
rect -515 -138 -513 -134
rect -509 -138 -507 -134
rect -515 -139 -507 -138
rect -505 -132 -497 -126
rect -505 -136 -503 -132
rect -499 -136 -497 -132
rect -505 -137 -497 -136
rect -495 -120 -488 -119
rect -495 -124 -493 -120
rect -489 -124 -488 -120
rect -495 -127 -488 -124
rect -495 -131 -493 -127
rect -489 -131 -488 -127
rect -284 -122 -283 -118
rect -279 -122 -277 -118
rect -284 -125 -277 -122
rect -284 -129 -283 -125
rect -279 -129 -277 -125
rect -284 -130 -277 -129
rect -495 -132 -488 -131
rect -495 -137 -490 -132
rect -282 -135 -277 -130
rect -275 -124 -269 -117
rect -191 -118 -184 -117
rect -191 -122 -190 -118
rect -186 -122 -184 -118
rect -275 -130 -267 -124
rect -275 -134 -273 -130
rect -269 -134 -267 -130
rect -275 -135 -267 -134
rect -505 -139 -499 -137
rect -273 -137 -267 -135
rect -265 -125 -257 -124
rect -265 -129 -263 -125
rect -259 -129 -257 -125
rect -265 -132 -257 -129
rect -265 -136 -263 -132
rect -259 -136 -257 -132
rect -265 -137 -257 -136
rect -255 -132 -248 -124
rect -191 -125 -184 -122
rect -191 -129 -190 -125
rect -186 -129 -184 -125
rect -191 -130 -184 -129
rect -255 -136 -253 -132
rect -249 -136 -248 -132
rect -189 -135 -184 -130
rect -182 -124 -176 -117
rect -104 -118 -97 -117
rect -104 -122 -103 -118
rect -99 -122 -97 -118
rect -182 -130 -174 -124
rect -182 -134 -180 -130
rect -176 -134 -174 -130
rect -182 -135 -174 -134
rect -255 -137 -248 -136
rect -180 -137 -174 -135
rect -172 -125 -164 -124
rect -172 -129 -170 -125
rect -166 -129 -164 -125
rect -172 -132 -164 -129
rect -172 -136 -170 -132
rect -166 -136 -164 -132
rect -172 -137 -164 -136
rect -162 -132 -155 -124
rect -104 -125 -97 -122
rect -104 -129 -103 -125
rect -99 -129 -97 -125
rect -104 -130 -97 -129
rect -162 -136 -160 -132
rect -156 -136 -155 -132
rect -102 -135 -97 -130
rect -95 -124 -89 -117
rect -95 -130 -87 -124
rect -95 -134 -93 -130
rect -89 -134 -87 -130
rect -95 -135 -87 -134
rect -162 -137 -155 -136
rect -93 -137 -87 -135
rect -85 -125 -77 -124
rect -85 -129 -83 -125
rect -79 -129 -77 -125
rect -85 -132 -77 -129
rect -85 -136 -83 -132
rect -79 -136 -77 -132
rect -85 -137 -77 -136
rect -75 -132 -68 -124
rect -75 -136 -73 -132
rect -69 -136 -68 -132
rect -17 -129 -2 -128
rect -13 -133 -2 -129
rect -17 -134 -2 -133
rect 0 -129 20 -128
rect 0 -133 16 -129
rect 0 -134 20 -133
rect 27 -129 37 -128
rect 27 -133 29 -129
rect 33 -133 37 -129
rect 27 -134 37 -133
rect 39 -129 58 -128
rect 39 -133 46 -129
rect 50 -133 58 -129
rect 39 -134 58 -133
rect 60 -129 68 -128
rect 60 -133 63 -129
rect 67 -133 68 -129
rect 60 -134 68 -133
rect 81 -129 91 -128
rect 81 -133 83 -129
rect 87 -133 91 -129
rect 81 -134 91 -133
rect 93 -129 112 -128
rect 93 -133 100 -129
rect 104 -133 112 -129
rect 93 -134 112 -133
rect 114 -129 122 -128
rect 114 -133 117 -129
rect 121 -133 122 -129
rect 114 -134 122 -133
rect 137 -129 147 -128
rect 137 -133 139 -129
rect 143 -133 147 -129
rect 137 -134 147 -133
rect 149 -129 168 -128
rect 149 -133 156 -129
rect 160 -133 168 -129
rect 149 -134 168 -133
rect 170 -129 178 -128
rect 170 -133 173 -129
rect 177 -133 178 -129
rect 170 -134 178 -133
rect 191 -129 201 -128
rect 191 -133 193 -129
rect 197 -133 201 -129
rect 191 -134 201 -133
rect 203 -129 222 -128
rect 203 -133 210 -129
rect 214 -133 222 -129
rect 203 -134 222 -133
rect 224 -129 232 -128
rect 224 -133 227 -129
rect 231 -133 232 -129
rect 224 -134 232 -133
rect -75 -137 -68 -136
rect -780 -187 -775 -181
rect -782 -188 -775 -187
rect -782 -192 -781 -188
rect -777 -192 -775 -188
rect -782 -193 -775 -192
rect -773 -183 -767 -181
rect -773 -188 -765 -183
rect -773 -192 -771 -188
rect -767 -192 -765 -188
rect -773 -193 -765 -192
rect -763 -188 -755 -183
rect -763 -192 -761 -188
rect -757 -192 -755 -188
rect -763 -193 -755 -192
rect -753 -184 -746 -183
rect -753 -188 -751 -184
rect -747 -188 -746 -184
rect -694 -186 -689 -165
rect -753 -193 -746 -188
rect -696 -187 -689 -186
rect -696 -191 -695 -187
rect -691 -191 -689 -187
rect -696 -192 -689 -191
rect -687 -166 -675 -165
rect -687 -170 -685 -166
rect -681 -170 -675 -166
rect -687 -173 -675 -170
rect -687 -177 -685 -173
rect -681 -174 -675 -173
rect -658 -174 -653 -165
rect -681 -177 -673 -174
rect -687 -192 -673 -177
rect -671 -187 -663 -174
rect -671 -191 -669 -187
rect -665 -191 -663 -187
rect -671 -192 -663 -191
rect -661 -180 -653 -174
rect -661 -184 -659 -180
rect -655 -184 -653 -180
rect -661 -192 -653 -184
rect -651 -171 -646 -165
rect -651 -172 -644 -171
rect -651 -176 -649 -172
rect -645 -176 -644 -172
rect -651 -177 -644 -176
rect -651 -192 -646 -177
rect -610 -186 -605 -165
rect -612 -187 -605 -186
rect -612 -191 -611 -187
rect -607 -191 -605 -187
rect -612 -192 -605 -191
rect -603 -166 -591 -165
rect -603 -170 -601 -166
rect -597 -170 -591 -166
rect -603 -173 -591 -170
rect -603 -177 -601 -173
rect -597 -174 -591 -173
rect -574 -174 -569 -165
rect -597 -177 -589 -174
rect -603 -192 -589 -177
rect -587 -187 -579 -174
rect -587 -191 -585 -187
rect -581 -191 -579 -187
rect -587 -192 -579 -191
rect -577 -180 -569 -174
rect -577 -184 -575 -180
rect -571 -184 -569 -180
rect -577 -192 -569 -184
rect -567 -171 -562 -165
rect -567 -172 -560 -171
rect -567 -176 -565 -172
rect -561 -176 -560 -172
rect -567 -177 -560 -176
rect -567 -192 -562 -177
rect -548 -187 -543 -181
rect -550 -188 -543 -187
rect -550 -192 -549 -188
rect -545 -192 -543 -188
rect -550 -193 -543 -192
rect -541 -183 -535 -181
rect -541 -188 -533 -183
rect -541 -192 -539 -188
rect -535 -192 -533 -188
rect -541 -193 -533 -192
rect -531 -188 -523 -183
rect -531 -192 -529 -188
rect -525 -192 -523 -188
rect -531 -193 -523 -192
rect -521 -184 -514 -183
rect -521 -188 -519 -184
rect -515 -188 -514 -184
rect -451 -185 -446 -179
rect -521 -193 -514 -188
rect -453 -186 -446 -185
rect -453 -190 -452 -186
rect -448 -190 -446 -186
rect -453 -191 -446 -190
rect -444 -181 -438 -179
rect -444 -186 -436 -181
rect -444 -190 -442 -186
rect -438 -190 -436 -186
rect -444 -191 -436 -190
rect -434 -186 -426 -181
rect -434 -190 -432 -186
rect -428 -190 -426 -186
rect -434 -191 -426 -190
rect -424 -182 -417 -181
rect -424 -186 -422 -182
rect -418 -186 -417 -182
rect -365 -184 -360 -163
rect -424 -191 -417 -186
rect -367 -185 -360 -184
rect -367 -189 -366 -185
rect -362 -189 -360 -185
rect -367 -190 -360 -189
rect -358 -164 -346 -163
rect -358 -168 -356 -164
rect -352 -168 -346 -164
rect -358 -171 -346 -168
rect -358 -175 -356 -171
rect -352 -172 -346 -171
rect -329 -172 -324 -163
rect -352 -175 -344 -172
rect -358 -190 -344 -175
rect -342 -185 -334 -172
rect -342 -189 -340 -185
rect -336 -189 -334 -185
rect -342 -190 -334 -189
rect -332 -178 -324 -172
rect -332 -182 -330 -178
rect -326 -182 -324 -178
rect -332 -190 -324 -182
rect -322 -169 -317 -163
rect -322 -170 -315 -169
rect -322 -174 -320 -170
rect -316 -174 -315 -170
rect -322 -175 -315 -174
rect -322 -190 -317 -175
rect -281 -184 -276 -163
rect -283 -185 -276 -184
rect -283 -189 -282 -185
rect -278 -189 -276 -185
rect -283 -190 -276 -189
rect -274 -164 -262 -163
rect -274 -168 -272 -164
rect -268 -168 -262 -164
rect -274 -171 -262 -168
rect -274 -175 -272 -171
rect -268 -172 -262 -171
rect -245 -172 -240 -163
rect -268 -175 -260 -172
rect -274 -190 -260 -175
rect -258 -185 -250 -172
rect -258 -189 -256 -185
rect -252 -189 -250 -185
rect -258 -190 -250 -189
rect -248 -178 -240 -172
rect -248 -182 -246 -178
rect -242 -182 -240 -178
rect -248 -190 -240 -182
rect -238 -169 -233 -163
rect -238 -170 -231 -169
rect -238 -174 -236 -170
rect -232 -174 -231 -170
rect -238 -175 -231 -174
rect -238 -190 -233 -175
rect -219 -185 -214 -179
rect -221 -186 -214 -185
rect -221 -190 -220 -186
rect -216 -190 -214 -186
rect -221 -191 -214 -190
rect -212 -181 -206 -179
rect -212 -186 -204 -181
rect -212 -190 -210 -186
rect -206 -190 -204 -186
rect -212 -191 -204 -190
rect -202 -186 -194 -181
rect -202 -190 -200 -186
rect -196 -190 -194 -186
rect -202 -191 -194 -190
rect -192 -182 -185 -181
rect -124 -182 -119 -176
rect -192 -186 -190 -182
rect -186 -186 -185 -182
rect -192 -191 -185 -186
rect -126 -183 -119 -182
rect -126 -187 -125 -183
rect -121 -187 -119 -183
rect -126 -188 -119 -187
rect -117 -178 -111 -176
rect -117 -183 -109 -178
rect -117 -187 -115 -183
rect -111 -187 -109 -183
rect -117 -188 -109 -187
rect -107 -183 -99 -178
rect -107 -187 -105 -183
rect -101 -187 -99 -183
rect -107 -188 -99 -187
rect -97 -179 -90 -178
rect -97 -183 -95 -179
rect -91 -183 -90 -179
rect -38 -181 -33 -160
rect -97 -188 -90 -183
rect -40 -182 -33 -181
rect -40 -186 -39 -182
rect -35 -186 -33 -182
rect -40 -187 -33 -186
rect -31 -161 -19 -160
rect -31 -165 -29 -161
rect -25 -165 -19 -161
rect -31 -168 -19 -165
rect -31 -172 -29 -168
rect -25 -169 -19 -168
rect -2 -169 3 -160
rect -25 -172 -17 -169
rect -31 -187 -17 -172
rect -15 -182 -7 -169
rect -15 -186 -13 -182
rect -9 -186 -7 -182
rect -15 -187 -7 -186
rect -5 -175 3 -169
rect -5 -179 -3 -175
rect 1 -179 3 -175
rect -5 -187 3 -179
rect 5 -166 10 -160
rect 5 -167 12 -166
rect 5 -171 7 -167
rect 11 -171 12 -167
rect 5 -172 12 -171
rect 5 -187 10 -172
rect 46 -181 51 -160
rect 44 -182 51 -181
rect 44 -186 45 -182
rect 49 -186 51 -182
rect 44 -187 51 -186
rect 53 -161 65 -160
rect 53 -165 55 -161
rect 59 -165 65 -161
rect 53 -168 65 -165
rect 53 -172 55 -168
rect 59 -169 65 -168
rect 82 -169 87 -160
rect 59 -172 67 -169
rect 53 -187 67 -172
rect 69 -182 77 -169
rect 69 -186 71 -182
rect 75 -186 77 -182
rect 69 -187 77 -186
rect 79 -175 87 -169
rect 79 -179 81 -175
rect 85 -179 87 -175
rect 79 -187 87 -179
rect 89 -166 94 -160
rect 89 -167 96 -166
rect 89 -171 91 -167
rect 95 -171 96 -167
rect 89 -172 96 -171
rect 89 -187 94 -172
rect 108 -182 113 -176
rect 106 -183 113 -182
rect 106 -187 107 -183
rect 111 -187 113 -183
rect 106 -188 113 -187
rect 115 -178 121 -176
rect 115 -183 123 -178
rect 115 -187 117 -183
rect 121 -187 123 -183
rect 115 -188 123 -187
rect 125 -183 133 -178
rect 125 -187 127 -183
rect 131 -187 133 -183
rect 125 -188 133 -187
rect 135 -179 142 -178
rect 135 -183 137 -179
rect 141 -183 142 -179
rect 135 -188 142 -183
rect -670 -277 -662 -274
rect -687 -282 -682 -277
rect -689 -283 -682 -282
rect -689 -287 -688 -283
rect -684 -287 -682 -283
rect -689 -288 -682 -287
rect -687 -295 -682 -288
rect -680 -295 -675 -277
rect -673 -286 -662 -277
rect -660 -280 -655 -274
rect -14 -272 -6 -269
rect -341 -275 -333 -272
rect -358 -280 -353 -275
rect -660 -281 -653 -280
rect -660 -285 -658 -281
rect -654 -285 -653 -281
rect -660 -286 -653 -285
rect -360 -281 -353 -280
rect -360 -285 -359 -281
rect -355 -285 -353 -281
rect -360 -286 -353 -285
rect -673 -290 -664 -286
rect -673 -294 -670 -290
rect -666 -294 -664 -290
rect -673 -295 -664 -294
rect -358 -293 -353 -286
rect -351 -293 -346 -275
rect -344 -284 -333 -275
rect -331 -278 -326 -272
rect -31 -277 -26 -272
rect -33 -278 -26 -277
rect -331 -279 -324 -278
rect -331 -283 -329 -279
rect -325 -283 -324 -279
rect -33 -282 -32 -278
rect -28 -282 -26 -278
rect -33 -283 -26 -282
rect -331 -284 -324 -283
rect -344 -288 -335 -284
rect -344 -292 -341 -288
rect -337 -292 -335 -288
rect -31 -290 -26 -283
rect -24 -290 -19 -272
rect -17 -281 -6 -272
rect -4 -275 1 -269
rect -4 -276 3 -275
rect -4 -280 -2 -276
rect 2 -280 3 -276
rect -4 -281 3 -280
rect -17 -285 -8 -281
rect -17 -289 -14 -285
rect -10 -289 -8 -285
rect -17 -290 -8 -289
rect -344 -293 -335 -292
rect -781 -333 -776 -327
rect -783 -334 -776 -333
rect -783 -338 -782 -334
rect -778 -338 -776 -334
rect -783 -339 -776 -338
rect -774 -329 -768 -327
rect -774 -334 -766 -329
rect -774 -338 -772 -334
rect -768 -338 -766 -334
rect -774 -339 -766 -338
rect -764 -334 -756 -329
rect -764 -338 -762 -334
rect -758 -338 -756 -334
rect -764 -339 -756 -338
rect -754 -330 -747 -329
rect -754 -334 -752 -330
rect -748 -334 -747 -330
rect -695 -332 -690 -311
rect -754 -339 -747 -334
rect -697 -333 -690 -332
rect -697 -337 -696 -333
rect -692 -337 -690 -333
rect -697 -338 -690 -337
rect -688 -312 -676 -311
rect -688 -316 -686 -312
rect -682 -316 -676 -312
rect -688 -319 -676 -316
rect -688 -323 -686 -319
rect -682 -320 -676 -319
rect -659 -320 -654 -311
rect -682 -323 -674 -320
rect -688 -338 -674 -323
rect -672 -333 -664 -320
rect -672 -337 -670 -333
rect -666 -337 -664 -333
rect -672 -338 -664 -337
rect -662 -326 -654 -320
rect -662 -330 -660 -326
rect -656 -330 -654 -326
rect -662 -338 -654 -330
rect -652 -317 -647 -311
rect -652 -318 -645 -317
rect -652 -322 -650 -318
rect -646 -322 -645 -318
rect -652 -323 -645 -322
rect -652 -338 -647 -323
rect -611 -332 -606 -311
rect -613 -333 -606 -332
rect -613 -337 -612 -333
rect -608 -337 -606 -333
rect -613 -338 -606 -337
rect -604 -312 -592 -311
rect -604 -316 -602 -312
rect -598 -316 -592 -312
rect -604 -319 -592 -316
rect -604 -323 -602 -319
rect -598 -320 -592 -319
rect -575 -320 -570 -311
rect -598 -323 -590 -320
rect -604 -338 -590 -323
rect -588 -333 -580 -320
rect -588 -337 -586 -333
rect -582 -337 -580 -333
rect -588 -338 -580 -337
rect -578 -326 -570 -320
rect -578 -330 -576 -326
rect -572 -330 -570 -326
rect -578 -338 -570 -330
rect -568 -317 -563 -311
rect -568 -318 -561 -317
rect -568 -322 -566 -318
rect -562 -322 -561 -318
rect -568 -323 -561 -322
rect -568 -338 -563 -323
rect -549 -333 -544 -327
rect -551 -334 -544 -333
rect -551 -338 -550 -334
rect -546 -338 -544 -334
rect -551 -339 -544 -338
rect -542 -329 -536 -327
rect -542 -334 -534 -329
rect -542 -338 -540 -334
rect -536 -338 -534 -334
rect -542 -339 -534 -338
rect -532 -334 -524 -329
rect -532 -338 -530 -334
rect -526 -338 -524 -334
rect -532 -339 -524 -338
rect -522 -330 -515 -329
rect -522 -334 -520 -330
rect -516 -334 -515 -330
rect -452 -331 -447 -325
rect -522 -339 -515 -334
rect -454 -332 -447 -331
rect -454 -336 -453 -332
rect -449 -336 -447 -332
rect -454 -337 -447 -336
rect -445 -327 -439 -325
rect -445 -332 -437 -327
rect -445 -336 -443 -332
rect -439 -336 -437 -332
rect -445 -337 -437 -336
rect -435 -332 -427 -327
rect -435 -336 -433 -332
rect -429 -336 -427 -332
rect -435 -337 -427 -336
rect -425 -328 -418 -327
rect -425 -332 -423 -328
rect -419 -332 -418 -328
rect -366 -330 -361 -309
rect -425 -337 -418 -332
rect -368 -331 -361 -330
rect -368 -335 -367 -331
rect -363 -335 -361 -331
rect -368 -336 -361 -335
rect -359 -310 -347 -309
rect -359 -314 -357 -310
rect -353 -314 -347 -310
rect -359 -317 -347 -314
rect -359 -321 -357 -317
rect -353 -318 -347 -317
rect -330 -318 -325 -309
rect -353 -321 -345 -318
rect -359 -336 -345 -321
rect -343 -331 -335 -318
rect -343 -335 -341 -331
rect -337 -335 -335 -331
rect -343 -336 -335 -335
rect -333 -324 -325 -318
rect -333 -328 -331 -324
rect -327 -328 -325 -324
rect -333 -336 -325 -328
rect -323 -315 -318 -309
rect -323 -316 -316 -315
rect -323 -320 -321 -316
rect -317 -320 -316 -316
rect -323 -321 -316 -320
rect -323 -336 -318 -321
rect -282 -330 -277 -309
rect -284 -331 -277 -330
rect -284 -335 -283 -331
rect -279 -335 -277 -331
rect -284 -336 -277 -335
rect -275 -310 -263 -309
rect -275 -314 -273 -310
rect -269 -314 -263 -310
rect -275 -317 -263 -314
rect -275 -321 -273 -317
rect -269 -318 -263 -317
rect -246 -318 -241 -309
rect -269 -321 -261 -318
rect -275 -336 -261 -321
rect -259 -331 -251 -318
rect -259 -335 -257 -331
rect -253 -335 -251 -331
rect -259 -336 -251 -335
rect -249 -324 -241 -318
rect -249 -328 -247 -324
rect -243 -328 -241 -324
rect -249 -336 -241 -328
rect -239 -315 -234 -309
rect -239 -316 -232 -315
rect -239 -320 -237 -316
rect -233 -320 -232 -316
rect -239 -321 -232 -320
rect -239 -336 -234 -321
rect -220 -331 -215 -325
rect -222 -332 -215 -331
rect -222 -336 -221 -332
rect -217 -336 -215 -332
rect -222 -337 -215 -336
rect -213 -327 -207 -325
rect -213 -332 -205 -327
rect -213 -336 -211 -332
rect -207 -336 -205 -332
rect -213 -337 -205 -336
rect -203 -332 -195 -327
rect -203 -336 -201 -332
rect -197 -336 -195 -332
rect -203 -337 -195 -336
rect -193 -328 -186 -327
rect -125 -328 -120 -322
rect -193 -332 -191 -328
rect -187 -332 -186 -328
rect -193 -337 -186 -332
rect -127 -329 -120 -328
rect -127 -333 -126 -329
rect -122 -333 -120 -329
rect -127 -334 -120 -333
rect -118 -324 -112 -322
rect -118 -329 -110 -324
rect -118 -333 -116 -329
rect -112 -333 -110 -329
rect -118 -334 -110 -333
rect -108 -329 -100 -324
rect -108 -333 -106 -329
rect -102 -333 -100 -329
rect -108 -334 -100 -333
rect -98 -325 -91 -324
rect -98 -329 -96 -325
rect -92 -329 -91 -325
rect -39 -327 -34 -306
rect -98 -334 -91 -329
rect -41 -328 -34 -327
rect -41 -332 -40 -328
rect -36 -332 -34 -328
rect -41 -333 -34 -332
rect -32 -307 -20 -306
rect -32 -311 -30 -307
rect -26 -311 -20 -307
rect -32 -314 -20 -311
rect -32 -318 -30 -314
rect -26 -315 -20 -314
rect -3 -315 2 -306
rect -26 -318 -18 -315
rect -32 -333 -18 -318
rect -16 -328 -8 -315
rect -16 -332 -14 -328
rect -10 -332 -8 -328
rect -16 -333 -8 -332
rect -6 -321 2 -315
rect -6 -325 -4 -321
rect 0 -325 2 -321
rect -6 -333 2 -325
rect 4 -312 9 -306
rect 4 -313 11 -312
rect 4 -317 6 -313
rect 10 -317 11 -313
rect 4 -318 11 -317
rect 4 -333 9 -318
rect 45 -327 50 -306
rect 43 -328 50 -327
rect 43 -332 44 -328
rect 48 -332 50 -328
rect 43 -333 50 -332
rect 52 -307 64 -306
rect 52 -311 54 -307
rect 58 -311 64 -307
rect 52 -314 64 -311
rect 52 -318 54 -314
rect 58 -315 64 -314
rect 81 -315 86 -306
rect 58 -318 66 -315
rect 52 -333 66 -318
rect 68 -328 76 -315
rect 68 -332 70 -328
rect 74 -332 76 -328
rect 68 -333 76 -332
rect 78 -321 86 -315
rect 78 -325 80 -321
rect 84 -325 86 -321
rect 78 -333 86 -325
rect 88 -312 93 -306
rect 88 -313 95 -312
rect 88 -317 90 -313
rect 94 -317 95 -313
rect 88 -318 95 -317
rect 88 -333 93 -318
rect 107 -328 112 -322
rect 105 -329 112 -328
rect 105 -333 106 -329
rect 110 -333 112 -329
rect 105 -334 112 -333
rect 114 -324 120 -322
rect 114 -329 122 -324
rect 114 -333 116 -329
rect 120 -333 122 -329
rect 114 -334 122 -333
rect 124 -329 132 -324
rect 124 -333 126 -329
rect 130 -333 132 -329
rect 124 -334 132 -333
rect 134 -325 141 -324
rect 134 -329 136 -325
rect 140 -329 141 -325
rect 134 -334 141 -329
rect -671 -423 -663 -420
rect -688 -428 -683 -423
rect -690 -429 -683 -428
rect -690 -433 -689 -429
rect -685 -433 -683 -429
rect -690 -434 -683 -433
rect -688 -441 -683 -434
rect -681 -441 -676 -423
rect -674 -432 -663 -423
rect -661 -426 -656 -420
rect -15 -418 -7 -415
rect -342 -421 -334 -418
rect -359 -426 -354 -421
rect -661 -427 -654 -426
rect -661 -431 -659 -427
rect -655 -431 -654 -427
rect -661 -432 -654 -431
rect -361 -427 -354 -426
rect -361 -431 -360 -427
rect -356 -431 -354 -427
rect -361 -432 -354 -431
rect -674 -436 -665 -432
rect -674 -440 -671 -436
rect -667 -440 -665 -436
rect -674 -441 -665 -440
rect -359 -439 -354 -432
rect -352 -439 -347 -421
rect -345 -430 -334 -421
rect -332 -424 -327 -418
rect -32 -423 -27 -418
rect -34 -424 -27 -423
rect -332 -425 -325 -424
rect -332 -429 -330 -425
rect -326 -429 -325 -425
rect -34 -428 -33 -424
rect -29 -428 -27 -424
rect -34 -429 -27 -428
rect -332 -430 -325 -429
rect -345 -434 -336 -430
rect -345 -438 -342 -434
rect -338 -438 -336 -434
rect -32 -436 -27 -429
rect -25 -436 -20 -418
rect -18 -427 -7 -418
rect -5 -421 0 -415
rect -5 -422 2 -421
rect -5 -426 -3 -422
rect 1 -426 2 -422
rect -5 -427 2 -426
rect -18 -431 -9 -427
rect -18 -435 -15 -431
rect -11 -435 -9 -431
rect -18 -436 -9 -435
rect -345 -439 -336 -438
rect -478 -468 -472 -466
rect -487 -473 -482 -468
rect -489 -474 -482 -473
rect -489 -478 -488 -474
rect -484 -478 -482 -474
rect -489 -481 -482 -478
rect -489 -485 -488 -481
rect -484 -485 -482 -481
rect -489 -486 -482 -485
rect -480 -469 -472 -468
rect -480 -473 -478 -469
rect -474 -473 -472 -469
rect -480 -479 -472 -473
rect -470 -467 -462 -466
rect -470 -471 -468 -467
rect -464 -471 -462 -467
rect -470 -474 -462 -471
rect -470 -478 -468 -474
rect -464 -478 -462 -474
rect -470 -479 -462 -478
rect -460 -467 -453 -466
rect -460 -471 -458 -467
rect -454 -471 -453 -467
rect -385 -468 -379 -466
rect -460 -479 -453 -471
rect -394 -473 -389 -468
rect -396 -474 -389 -473
rect -396 -478 -395 -474
rect -391 -478 -389 -474
rect -480 -486 -474 -479
rect -396 -481 -389 -478
rect -396 -485 -395 -481
rect -391 -485 -389 -481
rect -396 -486 -389 -485
rect -387 -469 -379 -468
rect -387 -473 -385 -469
rect -381 -473 -379 -469
rect -387 -479 -379 -473
rect -377 -467 -369 -466
rect -377 -471 -375 -467
rect -371 -471 -369 -467
rect -377 -474 -369 -471
rect -377 -478 -375 -474
rect -371 -478 -369 -474
rect -377 -479 -369 -478
rect -367 -467 -360 -466
rect -367 -471 -365 -467
rect -361 -471 -360 -467
rect -298 -468 -292 -466
rect -367 -479 -360 -471
rect -307 -473 -302 -468
rect -309 -474 -302 -473
rect -309 -478 -308 -474
rect -304 -478 -302 -474
rect -387 -486 -381 -479
rect -309 -481 -302 -478
rect -309 -485 -308 -481
rect -304 -485 -302 -481
rect -309 -486 -302 -485
rect -300 -469 -292 -468
rect -300 -473 -298 -469
rect -294 -473 -292 -469
rect -300 -479 -292 -473
rect -290 -467 -282 -466
rect -290 -471 -288 -467
rect -284 -471 -282 -467
rect -290 -474 -282 -471
rect -290 -478 -288 -474
rect -284 -478 -282 -474
rect -290 -479 -282 -478
rect -280 -467 -273 -466
rect -280 -471 -278 -467
rect -274 -471 -273 -467
rect -280 -479 -273 -471
rect -300 -486 -294 -479
<< metal1 >>
rect -120 -11 246 -8
rect -104 -30 -101 -11
rect -59 -28 -55 -26
rect -21 -30 -18 -11
rect 42 -30 45 -11
rect 52 -16 55 -11
rect 96 -30 99 -11
rect 106 -16 109 -11
rect 152 -30 155 -11
rect 162 -16 165 -11
rect 206 -30 209 -11
rect 216 -16 219 -11
rect -59 -45 -55 -34
rect -76 -49 -73 -46
rect -59 -55 -56 -45
rect -4 -50 -1 -47
rect -59 -59 -58 -55
rect 13 -56 16 -34
rect 26 -39 29 -34
rect 59 -39 62 -34
rect 26 -42 62 -39
rect 28 -50 30 -47
rect 50 -50 51 -47
rect 59 -51 62 -42
rect 80 -39 83 -34
rect 113 -39 116 -34
rect 80 -42 116 -39
rect 136 -39 139 -34
rect 169 -39 172 -34
rect 136 -42 172 -39
rect 190 -39 193 -34
rect 223 -39 226 -34
rect 190 -42 226 -39
rect 66 -51 69 -42
rect 80 -47 87 -46
rect 80 -49 84 -47
rect 101 -51 105 -48
rect 59 -54 69 -51
rect -785 -71 -344 -67
rect -785 -93 -781 -71
rect -59 -67 -56 -59
rect 13 -60 14 -56
rect 13 -68 16 -60
rect 59 -67 62 -54
rect 101 -55 104 -51
rect 113 -54 116 -42
rect 169 -43 172 -42
rect 137 -50 140 -47
rect 113 -57 132 -54
rect 113 -67 116 -57
rect 161 -53 164 -51
rect 149 -61 152 -55
rect 163 -57 164 -53
rect 161 -58 164 -57
rect 126 -64 152 -61
rect 169 -67 172 -47
rect 193 -51 194 -48
rect 212 -47 218 -46
rect 212 -49 215 -47
rect 193 -60 196 -51
rect 223 -52 226 -42
rect 195 -64 196 -60
rect 223 -67 226 -56
rect -93 -77 -90 -71
rect -21 -77 -18 -72
rect 25 -77 28 -71
rect 79 -77 82 -71
rect 135 -77 138 -71
rect 189 -77 192 -71
rect -703 -80 -702 -77
rect -487 -80 -294 -79
rect -288 -80 -244 -78
rect -703 -81 -244 -80
rect -195 -81 -151 -78
rect -117 -80 228 -77
rect -117 -81 -56 -80
rect -708 -82 -56 -81
rect -708 -84 -282 -82
rect -708 -88 -684 -84
rect -680 -88 -674 -84
rect -670 -88 -597 -84
rect -593 -88 -587 -84
rect -583 -88 -504 -84
rect -500 -88 -494 -84
rect -490 -85 -282 -84
rect -490 -88 -484 -85
rect -288 -86 -282 -85
rect -278 -86 -272 -82
rect -268 -85 -189 -82
rect -268 -86 -244 -85
rect -195 -86 -189 -85
rect -185 -86 -179 -82
rect -175 -85 -102 -82
rect -175 -86 -151 -85
rect -108 -86 -102 -85
rect -98 -86 -92 -82
rect -88 -85 -56 -82
rect 51 -83 56 -80
rect 157 -83 161 -80
rect -88 -86 -64 -85
rect -17 -86 232 -83
rect -17 -91 -14 -86
rect -704 -98 -703 -94
rect -699 -98 -684 -94
rect -704 -105 -692 -101
rect -697 -110 -692 -105
rect -688 -102 -684 -98
rect -680 -96 -668 -93
rect -680 -99 -673 -96
rect -669 -100 -668 -96
rect -617 -98 -616 -94
rect -612 -98 -597 -94
rect -673 -101 -668 -100
rect -688 -106 -676 -102
rect -680 -110 -676 -106
rect -697 -114 -690 -110
rect -686 -114 -683 -110
rect -704 -127 -700 -118
rect -696 -122 -691 -118
rect -680 -125 -676 -114
rect -672 -115 -668 -101
rect -616 -105 -605 -101
rect -610 -110 -605 -105
rect -601 -102 -597 -98
rect -593 -96 -581 -93
rect -593 -99 -586 -96
rect -582 -100 -581 -96
rect -524 -98 -523 -94
rect -519 -98 -504 -94
rect -586 -101 -581 -100
rect -601 -106 -589 -102
rect -593 -110 -589 -106
rect -610 -114 -603 -110
rect -599 -114 -596 -110
rect -672 -118 -643 -115
rect -672 -119 -668 -118
rect -711 -131 -700 -127
rect -693 -127 -676 -125
rect -689 -129 -676 -127
rect -673 -120 -668 -119
rect -669 -124 -668 -120
rect -673 -127 -668 -124
rect -693 -134 -689 -131
rect -669 -131 -668 -127
rect -673 -132 -668 -131
rect -704 -138 -703 -134
rect -699 -138 -698 -134
rect -704 -144 -698 -138
rect -693 -139 -689 -138
rect -684 -136 -683 -132
rect -679 -136 -678 -132
rect -684 -144 -678 -136
rect -708 -148 -674 -144
rect -670 -148 -664 -144
rect -708 -152 -664 -148
rect -707 -159 -703 -152
rect -647 -154 -643 -118
rect -617 -128 -613 -118
rect -609 -122 -604 -118
rect -593 -125 -589 -114
rect -585 -119 -581 -101
rect -523 -105 -512 -101
rect -517 -110 -512 -105
rect -508 -102 -504 -98
rect -500 -96 -488 -93
rect -284 -94 -272 -91
rect -500 -99 -493 -96
rect -489 -100 -488 -96
rect -475 -100 -303 -96
rect -298 -100 -297 -96
rect -284 -98 -283 -94
rect -279 -97 -272 -94
rect -268 -96 -253 -92
rect -249 -96 -248 -92
rect -191 -94 -179 -91
rect -284 -99 -279 -98
rect -493 -101 -488 -100
rect -508 -106 -496 -102
rect -500 -110 -496 -106
rect -517 -114 -510 -110
rect -506 -114 -503 -110
rect -620 -131 -613 -128
rect -606 -127 -589 -125
rect -602 -129 -589 -127
rect -586 -120 -581 -119
rect -582 -124 -581 -120
rect -586 -127 -581 -124
rect -606 -134 -602 -131
rect -582 -129 -581 -127
rect -582 -131 -575 -129
rect -586 -132 -575 -131
rect -524 -128 -520 -118
rect -516 -122 -511 -118
rect -500 -125 -496 -114
rect -492 -119 -488 -101
rect -284 -106 -280 -99
rect -268 -100 -264 -96
rect -191 -98 -190 -94
rect -186 -97 -179 -94
rect -175 -96 -160 -92
rect -156 -96 -155 -92
rect -104 -94 -92 -91
rect -191 -99 -186 -98
rect -340 -110 -280 -106
rect -284 -117 -280 -110
rect -276 -104 -264 -100
rect -260 -102 -249 -99
rect -276 -108 -272 -104
rect -260 -108 -255 -102
rect -269 -112 -266 -108
rect -262 -112 -255 -108
rect -191 -110 -187 -99
rect -175 -100 -171 -96
rect -104 -98 -103 -94
rect -99 -97 -92 -94
rect -88 -96 -73 -92
rect -69 -96 -68 -92
rect 29 -92 32 -86
rect 83 -92 86 -86
rect 139 -92 142 -86
rect 193 -92 196 -86
rect -104 -99 -99 -98
rect -284 -118 -279 -117
rect -527 -131 -520 -128
rect -513 -127 -496 -125
rect -509 -129 -496 -127
rect -493 -120 -488 -119
rect -489 -124 -488 -120
rect -475 -122 -302 -119
rect -284 -122 -283 -118
rect -493 -127 -488 -124
rect -617 -138 -616 -134
rect -612 -138 -611 -134
rect -617 -144 -611 -138
rect -606 -139 -602 -138
rect -597 -136 -596 -132
rect -592 -136 -591 -132
rect -513 -134 -509 -131
rect -489 -131 -488 -127
rect -284 -125 -279 -122
rect -284 -129 -283 -125
rect -276 -123 -272 -112
rect -214 -113 -187 -110
rect -261 -120 -256 -116
rect -276 -125 -259 -123
rect -276 -127 -263 -125
rect -284 -130 -279 -129
rect -252 -126 -248 -116
rect -214 -125 -210 -113
rect -252 -129 -245 -126
rect -493 -132 -488 -131
rect -597 -144 -591 -136
rect -524 -138 -523 -134
rect -519 -138 -518 -134
rect -524 -144 -518 -138
rect -513 -139 -509 -138
rect -504 -136 -503 -132
rect -499 -136 -498 -132
rect -274 -134 -273 -130
rect -269 -134 -268 -130
rect -504 -144 -498 -136
rect -475 -140 -301 -137
rect -274 -142 -268 -134
rect -263 -132 -259 -129
rect -191 -117 -187 -113
rect -183 -104 -171 -100
rect -167 -100 -153 -99
rect -167 -102 -156 -100
rect -183 -108 -179 -104
rect -167 -108 -162 -102
rect -176 -112 -173 -108
rect -169 -112 -162 -108
rect -191 -118 -186 -117
rect -191 -122 -190 -118
rect -191 -125 -186 -122
rect -191 -129 -190 -125
rect -183 -123 -179 -112
rect -104 -113 -100 -99
rect -88 -100 -84 -96
rect -168 -120 -163 -116
rect -183 -125 -166 -123
rect -183 -127 -170 -125
rect -191 -130 -186 -129
rect -159 -126 -155 -116
rect -126 -117 -100 -113
rect -96 -104 -84 -100
rect -80 -100 -66 -99
rect -80 -102 -69 -100
rect -96 -108 -92 -104
rect -80 -108 -75 -102
rect -41 -100 10 -99
rect -41 -102 14 -100
rect 17 -103 20 -95
rect -89 -112 -86 -108
rect -82 -112 -75 -108
rect 17 -107 18 -103
rect -159 -129 -152 -126
rect -140 -127 -139 -123
rect -263 -137 -259 -136
rect -254 -136 -253 -132
rect -249 -136 -248 -132
rect -254 -142 -248 -136
rect -181 -134 -180 -130
rect -176 -134 -175 -130
rect -181 -142 -175 -134
rect -170 -132 -166 -129
rect -170 -137 -166 -136
rect -161 -136 -160 -132
rect -156 -136 -155 -132
rect -161 -142 -155 -136
rect -621 -148 -587 -144
rect -583 -148 -577 -144
rect -621 -149 -577 -148
rect -528 -148 -494 -144
rect -490 -148 -484 -144
rect -621 -152 -594 -149
rect -528 -152 -484 -148
rect -288 -146 -282 -142
rect -278 -146 -244 -142
rect -195 -146 -189 -142
rect -185 -146 -151 -142
rect -288 -150 -244 -146
rect -619 -159 -615 -152
rect -582 -156 -549 -153
rect -528 -159 -524 -152
rect -252 -154 -248 -150
rect -233 -151 -203 -148
rect -195 -150 -151 -146
rect -140 -147 -136 -127
rect -294 -155 -190 -154
rect -294 -157 -168 -155
rect -159 -157 -155 -150
rect -126 -148 -122 -117
rect -104 -118 -99 -117
rect -104 -122 -103 -118
rect -116 -147 -112 -127
rect -104 -125 -99 -122
rect -104 -129 -103 -125
rect -96 -123 -92 -112
rect 0 -116 3 -113
rect -81 -120 -76 -116
rect -96 -125 -79 -123
rect -96 -127 -83 -125
rect -104 -130 -99 -129
rect -72 -125 -68 -116
rect -72 -129 -64 -125
rect 17 -129 20 -107
rect 63 -109 66 -96
rect 78 -100 100 -99
rect 74 -102 100 -100
rect 63 -112 72 -109
rect 32 -116 34 -113
rect 54 -116 55 -113
rect 30 -121 33 -120
rect 63 -121 66 -112
rect 69 -118 72 -112
rect 84 -116 88 -114
rect 97 -113 100 -102
rect 84 -117 91 -116
rect 105 -112 108 -108
rect 117 -106 120 -96
rect 117 -109 136 -106
rect 165 -106 168 -105
rect 105 -115 109 -112
rect 69 -121 76 -118
rect 30 -124 66 -121
rect 30 -129 33 -124
rect 63 -129 66 -124
rect 117 -123 120 -109
rect 167 -110 168 -106
rect 165 -112 168 -110
rect 141 -116 144 -113
rect 173 -116 176 -96
rect 199 -103 200 -99
rect 197 -112 200 -103
rect 227 -107 230 -96
rect 197 -115 198 -112
rect 216 -116 219 -114
rect 216 -117 222 -116
rect 173 -121 176 -120
rect 227 -121 230 -111
rect 84 -126 120 -123
rect 84 -129 87 -126
rect 117 -129 120 -126
rect 140 -124 176 -121
rect 140 -129 143 -124
rect 173 -129 176 -124
rect 194 -124 230 -121
rect 194 -129 197 -124
rect 227 -129 230 -124
rect -94 -134 -93 -130
rect -89 -134 -88 -130
rect -94 -142 -88 -134
rect -83 -132 -79 -129
rect -83 -137 -79 -136
rect -74 -136 -73 -132
rect -69 -136 -68 -132
rect -74 -142 -68 -136
rect -108 -146 -102 -142
rect -98 -146 -64 -142
rect -108 -150 -64 -146
rect -70 -157 -66 -150
rect -17 -152 -14 -133
rect 46 -152 49 -133
rect 56 -152 59 -147
rect 100 -152 103 -133
rect 110 -152 113 -147
rect 156 -152 159 -133
rect 166 -152 169 -147
rect 210 -152 213 -133
rect 220 -152 223 -147
rect 241 -152 246 -11
rect -19 -154 246 -152
rect -56 -155 246 -154
rect -56 -157 146 -155
rect -512 -158 146 -157
rect -512 -159 -124 -158
rect -816 -160 -589 -159
rect -576 -160 -124 -159
rect -816 -161 -124 -160
rect -816 -163 -451 -161
rect -816 -167 -780 -163
rect -776 -167 -766 -163
rect -762 -167 -752 -163
rect -748 -166 -669 -163
rect -748 -167 -685 -166
rect -816 -278 -812 -167
rect -796 -168 -781 -167
rect -782 -187 -778 -180
rect -782 -188 -777 -187
rect -782 -192 -781 -188
rect -774 -188 -770 -167
rect -767 -173 -754 -172
rect -767 -177 -764 -173
rect -760 -177 -758 -173
rect -767 -178 -754 -177
rect -767 -185 -761 -178
rect -751 -184 -747 -167
rect -681 -167 -669 -166
rect -665 -166 -585 -163
rect -665 -167 -601 -166
rect -704 -178 -692 -172
rect -685 -173 -681 -170
rect -597 -167 -585 -166
rect -581 -167 -548 -163
rect -544 -167 -534 -163
rect -530 -167 -520 -163
rect -516 -165 -451 -163
rect -447 -165 -437 -161
rect -433 -165 -423 -161
rect -419 -164 -340 -161
rect -419 -165 -356 -164
rect -516 -167 -481 -165
rect -671 -176 -649 -172
rect -645 -176 -644 -172
rect -620 -173 -608 -172
rect -671 -177 -667 -176
rect -685 -178 -681 -177
rect -704 -181 -699 -178
rect -704 -182 -703 -181
rect -774 -192 -771 -188
rect -767 -192 -766 -188
rect -762 -192 -761 -188
rect -757 -192 -756 -188
rect -751 -189 -747 -188
rect -712 -185 -703 -182
rect -678 -181 -667 -177
rect -620 -177 -615 -173
rect -611 -177 -608 -173
rect -620 -178 -608 -177
rect -601 -173 -597 -170
rect -587 -176 -565 -172
rect -561 -176 -560 -172
rect -587 -177 -583 -176
rect -601 -178 -597 -177
rect -678 -185 -674 -181
rect -660 -184 -659 -180
rect -655 -184 -644 -180
rect -782 -193 -777 -192
rect -782 -201 -778 -193
rect -762 -197 -756 -192
rect -775 -201 -774 -197
rect -770 -201 -756 -197
rect -750 -199 -746 -196
rect -712 -199 -709 -185
rect -704 -186 -699 -185
rect -695 -187 -674 -185
rect -782 -210 -778 -205
rect -782 -211 -777 -210
rect -782 -215 -781 -211
rect -777 -215 -770 -212
rect -782 -218 -770 -215
rect -766 -214 -762 -201
rect -703 -191 -695 -190
rect -691 -189 -674 -187
rect -703 -194 -691 -191
rect -750 -205 -746 -203
rect -759 -209 -755 -205
rect -751 -209 -746 -205
rect -759 -210 -746 -209
rect -703 -206 -699 -194
rect -678 -196 -674 -189
rect -670 -191 -669 -187
rect -665 -188 -664 -187
rect -665 -191 -653 -188
rect -670 -192 -653 -191
rect -657 -195 -653 -192
rect -657 -196 -652 -195
rect -689 -202 -683 -197
rect -678 -200 -666 -196
rect -662 -200 -661 -196
rect -657 -200 -656 -196
rect -689 -204 -687 -202
rect -696 -206 -687 -204
rect -657 -201 -652 -200
rect -648 -200 -644 -184
rect -620 -181 -615 -178
rect -620 -185 -619 -181
rect -594 -181 -583 -177
rect -594 -185 -590 -181
rect -576 -184 -575 -180
rect -571 -184 -560 -180
rect -620 -186 -615 -185
rect -611 -187 -590 -185
rect -619 -191 -611 -190
rect -607 -189 -590 -187
rect -619 -194 -607 -191
rect -657 -205 -653 -201
rect -696 -210 -683 -206
rect -677 -209 -653 -205
rect -648 -204 -646 -200
rect -703 -211 -699 -210
rect -677 -211 -673 -209
rect -766 -218 -752 -214
rect -748 -218 -747 -214
rect -690 -218 -689 -214
rect -685 -218 -684 -214
rect -648 -213 -644 -204
rect -619 -206 -615 -194
rect -594 -196 -590 -189
rect -586 -191 -585 -187
rect -581 -188 -580 -187
rect -581 -191 -569 -188
rect -586 -192 -569 -191
rect -573 -195 -569 -192
rect -573 -196 -568 -195
rect -605 -202 -599 -197
rect -594 -200 -582 -196
rect -578 -200 -577 -196
rect -573 -200 -572 -196
rect -605 -204 -603 -202
rect -612 -206 -603 -204
rect -573 -201 -568 -200
rect -573 -205 -569 -201
rect -612 -210 -599 -206
rect -593 -209 -569 -205
rect -619 -211 -615 -210
rect -593 -211 -589 -209
rect -677 -216 -673 -215
rect -668 -217 -667 -213
rect -663 -217 -644 -213
rect -690 -223 -684 -218
rect -606 -218 -605 -214
rect -601 -218 -600 -214
rect -564 -213 -560 -184
rect -550 -187 -546 -180
rect -550 -188 -545 -187
rect -550 -192 -549 -188
rect -542 -188 -538 -167
rect -535 -173 -522 -172
rect -535 -177 -532 -173
rect -528 -177 -526 -173
rect -535 -178 -522 -177
rect -535 -185 -529 -178
rect -519 -184 -515 -167
rect -542 -192 -539 -188
rect -535 -192 -534 -188
rect -530 -192 -529 -188
rect -525 -192 -524 -188
rect -519 -189 -515 -188
rect -550 -193 -545 -192
rect -550 -201 -546 -193
rect -530 -197 -524 -192
rect -543 -201 -542 -197
rect -538 -201 -524 -197
rect -518 -198 -514 -196
rect -593 -216 -589 -215
rect -584 -217 -583 -213
rect -579 -217 -560 -213
rect -556 -204 -546 -201
rect -556 -216 -553 -204
rect -606 -223 -600 -218
rect -550 -210 -546 -204
rect -550 -211 -545 -210
rect -550 -215 -549 -211
rect -545 -215 -538 -212
rect -550 -218 -538 -215
rect -534 -214 -530 -201
rect -518 -205 -514 -202
rect -527 -209 -523 -205
rect -519 -209 -514 -205
rect -527 -210 -514 -209
rect -534 -218 -520 -214
rect -516 -218 -515 -214
rect -783 -227 -780 -223
rect -776 -227 -770 -223
rect -766 -227 -702 -223
rect -698 -227 -649 -223
rect -645 -227 -618 -223
rect -614 -227 -565 -223
rect -561 -227 -548 -223
rect -544 -227 -538 -223
rect -534 -224 -510 -223
rect -534 -227 -516 -224
rect -797 -230 -516 -227
rect -797 -231 -510 -230
rect -693 -233 -649 -231
rect -693 -237 -687 -233
rect -683 -237 -659 -233
rect -655 -237 -649 -233
rect -689 -245 -683 -237
rect -689 -249 -688 -245
rect -684 -249 -683 -245
rect -678 -245 -674 -244
rect -669 -245 -663 -237
rect -669 -249 -668 -245
rect -664 -249 -663 -245
rect -658 -245 -653 -242
rect -654 -249 -653 -245
rect -678 -252 -674 -249
rect -658 -250 -653 -249
rect -678 -256 -661 -252
rect -689 -268 -685 -258
rect -681 -263 -676 -259
rect -665 -260 -661 -256
rect -681 -271 -675 -267
rect -671 -271 -668 -267
rect -817 -298 -812 -278
rect -681 -277 -677 -271
rect -665 -275 -661 -264
rect -694 -280 -677 -277
rect -673 -279 -661 -275
rect -657 -254 -496 -250
rect -673 -283 -669 -279
rect -657 -280 -653 -254
rect -487 -276 -483 -167
rect -453 -185 -449 -178
rect -453 -186 -448 -185
rect -453 -190 -452 -186
rect -445 -186 -441 -165
rect -438 -171 -425 -170
rect -438 -175 -435 -171
rect -431 -175 -429 -171
rect -438 -176 -425 -175
rect -438 -183 -432 -176
rect -422 -182 -418 -165
rect -352 -165 -340 -164
rect -336 -164 -256 -161
rect -336 -165 -272 -164
rect -375 -176 -363 -170
rect -356 -171 -352 -168
rect -268 -165 -256 -164
rect -252 -165 -219 -161
rect -215 -165 -205 -161
rect -201 -165 -191 -161
rect -187 -162 -124 -161
rect -120 -162 -110 -158
rect -106 -162 -96 -158
rect -92 -161 -13 -158
rect -92 -162 -29 -161
rect -187 -165 -151 -162
rect -342 -174 -320 -170
rect -316 -174 -315 -170
rect -300 -171 -279 -170
rect -342 -175 -338 -174
rect -356 -176 -352 -175
rect -375 -179 -370 -176
rect -375 -180 -374 -179
rect -445 -190 -442 -186
rect -438 -190 -437 -186
rect -433 -190 -432 -186
rect -428 -190 -427 -186
rect -422 -187 -418 -186
rect -383 -183 -374 -180
rect -349 -179 -338 -175
rect -300 -175 -286 -171
rect -282 -175 -279 -171
rect -300 -176 -279 -175
rect -272 -171 -268 -168
rect -258 -174 -236 -170
rect -232 -174 -231 -170
rect -258 -175 -254 -174
rect -272 -176 -268 -175
rect -349 -183 -345 -179
rect -331 -182 -330 -178
rect -326 -182 -315 -178
rect -453 -191 -448 -190
rect -453 -199 -449 -191
rect -433 -195 -427 -190
rect -446 -199 -445 -195
rect -441 -199 -427 -195
rect -421 -197 -417 -194
rect -383 -197 -380 -183
rect -375 -184 -370 -183
rect -366 -185 -345 -183
rect -453 -208 -449 -203
rect -453 -209 -448 -208
rect -453 -213 -452 -209
rect -448 -213 -441 -210
rect -453 -216 -441 -213
rect -437 -212 -433 -199
rect -374 -189 -366 -188
rect -362 -187 -345 -185
rect -374 -192 -362 -189
rect -421 -203 -417 -201
rect -430 -207 -426 -203
rect -422 -207 -417 -203
rect -430 -208 -417 -207
rect -374 -204 -370 -192
rect -349 -194 -345 -187
rect -341 -189 -340 -185
rect -336 -186 -335 -185
rect -336 -189 -324 -186
rect -341 -190 -324 -189
rect -328 -193 -324 -190
rect -328 -194 -323 -193
rect -360 -200 -354 -195
rect -349 -198 -337 -194
rect -333 -198 -332 -194
rect -328 -198 -327 -194
rect -360 -202 -358 -200
rect -367 -204 -358 -202
rect -328 -199 -323 -198
rect -319 -198 -315 -182
rect -291 -179 -286 -176
rect -291 -183 -290 -179
rect -265 -179 -254 -175
rect -265 -183 -261 -179
rect -247 -182 -246 -178
rect -242 -182 -229 -178
rect -291 -184 -286 -183
rect -282 -185 -261 -183
rect -290 -189 -282 -188
rect -278 -187 -261 -185
rect -290 -192 -278 -189
rect -328 -203 -324 -199
rect -367 -208 -354 -204
rect -348 -207 -324 -203
rect -319 -202 -317 -198
rect -374 -209 -370 -208
rect -348 -209 -344 -207
rect -437 -216 -423 -212
rect -419 -216 -418 -212
rect -361 -216 -360 -212
rect -356 -216 -355 -212
rect -319 -211 -315 -202
rect -290 -204 -286 -192
rect -265 -194 -261 -187
rect -257 -189 -256 -185
rect -252 -186 -251 -185
rect -252 -189 -240 -186
rect -257 -190 -240 -189
rect -244 -193 -240 -190
rect -244 -194 -239 -193
rect -276 -200 -270 -195
rect -265 -198 -253 -194
rect -249 -198 -248 -194
rect -244 -198 -243 -194
rect -276 -202 -274 -200
rect -283 -204 -274 -202
rect -244 -199 -239 -198
rect -244 -203 -240 -199
rect -283 -208 -270 -204
rect -264 -207 -240 -203
rect -290 -209 -286 -208
rect -264 -209 -260 -207
rect -348 -214 -344 -213
rect -339 -215 -338 -211
rect -334 -215 -315 -211
rect -361 -221 -355 -216
rect -277 -216 -276 -212
rect -272 -216 -271 -212
rect -235 -211 -231 -182
rect -221 -185 -217 -178
rect -221 -186 -216 -185
rect -221 -190 -220 -186
rect -213 -186 -209 -165
rect -206 -171 -193 -170
rect -206 -175 -203 -171
rect -199 -175 -197 -171
rect -206 -176 -193 -175
rect -206 -183 -200 -176
rect -190 -182 -186 -165
rect -213 -190 -210 -186
rect -206 -190 -205 -186
rect -201 -190 -200 -186
rect -196 -190 -195 -186
rect -190 -187 -186 -186
rect -221 -191 -216 -190
rect -221 -199 -217 -191
rect -201 -195 -195 -190
rect -214 -199 -213 -195
rect -209 -199 -195 -195
rect -189 -196 -185 -194
rect -264 -214 -260 -213
rect -255 -215 -254 -211
rect -250 -215 -231 -211
rect -227 -202 -217 -199
rect -227 -214 -224 -202
rect -277 -221 -271 -216
rect -221 -208 -217 -202
rect -221 -209 -216 -208
rect -221 -213 -220 -209
rect -216 -213 -209 -210
rect -221 -216 -209 -213
rect -205 -212 -201 -199
rect -189 -203 -185 -200
rect -198 -207 -194 -203
rect -190 -207 -185 -203
rect -198 -208 -185 -207
rect -205 -216 -191 -212
rect -187 -216 -186 -212
rect -454 -225 -451 -221
rect -447 -225 -441 -221
rect -437 -225 -373 -221
rect -369 -225 -320 -221
rect -316 -225 -289 -221
rect -285 -225 -236 -221
rect -232 -225 -219 -221
rect -215 -225 -209 -221
rect -205 -222 -181 -221
rect -205 -225 -189 -222
rect -454 -226 -189 -225
rect -469 -228 -189 -226
rect -183 -228 -181 -222
rect -469 -229 -181 -228
rect -469 -230 -453 -229
rect -364 -231 -320 -229
rect -364 -235 -358 -231
rect -354 -235 -330 -231
rect -326 -235 -320 -231
rect -360 -243 -354 -235
rect -360 -247 -359 -243
rect -355 -247 -354 -243
rect -349 -243 -345 -242
rect -340 -243 -334 -235
rect -340 -247 -339 -243
rect -335 -247 -334 -243
rect -329 -243 -324 -240
rect -325 -247 -324 -243
rect -349 -250 -345 -247
rect -329 -248 -324 -247
rect -467 -254 -399 -250
rect -349 -254 -332 -250
rect -360 -266 -356 -256
rect -352 -261 -347 -257
rect -336 -258 -332 -254
rect -352 -269 -346 -265
rect -342 -269 -339 -265
rect -658 -281 -653 -280
rect -689 -287 -688 -283
rect -684 -287 -669 -283
rect -666 -285 -658 -283
rect -654 -285 -653 -281
rect -666 -287 -653 -285
rect -671 -293 -670 -290
rect -693 -294 -670 -293
rect -666 -293 -665 -290
rect -666 -294 -659 -293
rect -693 -297 -659 -294
rect -655 -297 -649 -293
rect -693 -298 -649 -297
rect -488 -296 -483 -276
rect -352 -275 -348 -269
rect -336 -273 -332 -262
rect -365 -278 -348 -275
rect -344 -277 -332 -273
rect -328 -254 -324 -248
rect -328 -257 -177 -254
rect -173 -257 -172 -254
rect -344 -281 -340 -277
rect -328 -278 -324 -257
rect -160 -273 -156 -165
rect -126 -182 -122 -175
rect -126 -183 -121 -182
rect -126 -187 -125 -183
rect -118 -183 -114 -162
rect -111 -168 -98 -167
rect -111 -172 -108 -168
rect -104 -172 -102 -168
rect -111 -173 -98 -172
rect -111 -180 -105 -173
rect -95 -179 -91 -162
rect -25 -162 -13 -161
rect -9 -161 71 -158
rect -9 -162 55 -161
rect -48 -173 -36 -167
rect -29 -168 -25 -165
rect 59 -162 71 -161
rect 75 -162 108 -158
rect 112 -162 122 -158
rect 126 -162 136 -158
rect 140 -162 146 -158
rect -15 -171 7 -167
rect 11 -171 12 -167
rect 25 -168 48 -167
rect -15 -172 -11 -171
rect 25 -172 41 -168
rect 45 -172 48 -168
rect -29 -173 -25 -172
rect -48 -176 -43 -173
rect -48 -177 -47 -176
rect -118 -187 -115 -183
rect -111 -187 -110 -183
rect -106 -187 -105 -183
rect -101 -187 -100 -183
rect -95 -184 -91 -183
rect -126 -188 -121 -187
rect -126 -196 -122 -188
rect -106 -192 -100 -187
rect -119 -196 -118 -192
rect -114 -196 -100 -192
rect -94 -194 -90 -191
rect -126 -205 -122 -200
rect -126 -206 -121 -205
rect -126 -210 -125 -206
rect -121 -210 -114 -207
rect -126 -213 -114 -210
rect -110 -209 -106 -196
rect -94 -200 -90 -198
rect -103 -204 -99 -200
rect -95 -204 -90 -200
rect -103 -205 -90 -204
rect -110 -213 -96 -209
rect -92 -213 -91 -209
rect -67 -211 -63 -182
rect -56 -180 -47 -177
rect -22 -176 -11 -172
rect -22 -180 -18 -176
rect -4 -179 -3 -175
rect 1 -179 12 -175
rect -56 -194 -53 -180
rect -48 -181 -43 -180
rect -39 -182 -18 -180
rect -47 -186 -39 -185
rect -35 -184 -18 -182
rect -47 -189 -35 -186
rect -47 -201 -43 -189
rect -22 -191 -18 -184
rect -14 -186 -13 -182
rect -9 -183 -8 -182
rect -9 -186 3 -183
rect -14 -187 3 -186
rect -1 -190 3 -187
rect -1 -191 4 -190
rect -33 -197 -27 -192
rect -22 -195 -10 -191
rect -6 -195 -5 -191
rect -1 -195 0 -191
rect -33 -199 -31 -197
rect -40 -201 -31 -199
rect -1 -196 4 -195
rect 8 -195 12 -179
rect -1 -200 3 -196
rect -40 -205 -27 -201
rect -21 -204 3 -200
rect 8 -199 10 -195
rect -47 -206 -43 -205
rect -21 -206 -17 -204
rect -67 -215 -66 -211
rect -34 -213 -33 -209
rect -29 -213 -28 -209
rect 8 -208 12 -199
rect -21 -211 -17 -210
rect -12 -212 -11 -208
rect -7 -212 12 -208
rect 19 -211 22 -180
rect -34 -218 -28 -213
rect 26 -218 30 -172
rect 36 -173 48 -172
rect 55 -168 59 -165
rect 69 -171 91 -167
rect 95 -171 96 -167
rect 69 -172 73 -171
rect 55 -173 59 -172
rect 36 -176 41 -173
rect 36 -180 37 -176
rect 62 -176 73 -172
rect 62 -180 66 -176
rect 80 -179 81 -175
rect 85 -179 96 -175
rect 36 -181 41 -180
rect 45 -182 66 -180
rect 37 -186 45 -185
rect 49 -184 66 -182
rect 37 -189 49 -186
rect 37 -201 41 -189
rect 62 -191 66 -184
rect 70 -186 71 -182
rect 75 -183 76 -182
rect 75 -186 87 -183
rect 70 -187 87 -186
rect 83 -190 87 -187
rect 83 -191 88 -190
rect 51 -197 57 -192
rect 62 -195 74 -191
rect 78 -195 79 -191
rect 83 -195 84 -191
rect 51 -199 53 -197
rect 44 -201 53 -199
rect 83 -196 88 -195
rect 83 -200 87 -196
rect 44 -205 57 -201
rect 63 -204 87 -200
rect 37 -206 41 -205
rect 63 -206 67 -204
rect 50 -213 51 -209
rect 55 -213 56 -209
rect 92 -208 96 -179
rect 106 -182 110 -175
rect 106 -183 111 -182
rect 106 -187 107 -183
rect 114 -183 118 -162
rect 121 -168 134 -167
rect 121 -172 124 -168
rect 128 -172 130 -168
rect 121 -173 134 -172
rect 121 -180 127 -173
rect 137 -179 141 -162
rect 114 -187 117 -183
rect 121 -187 122 -183
rect 126 -187 127 -183
rect 131 -187 132 -183
rect 137 -184 141 -183
rect 106 -188 111 -187
rect 106 -196 110 -188
rect 126 -192 132 -187
rect 113 -196 114 -192
rect 118 -196 132 -192
rect 138 -193 142 -191
rect 63 -211 67 -210
rect 72 -212 73 -208
rect 77 -212 96 -208
rect 100 -199 110 -196
rect 100 -211 103 -199
rect 50 -218 56 -213
rect 106 -205 110 -199
rect 106 -206 111 -205
rect 106 -210 107 -206
rect 111 -210 118 -207
rect 106 -213 118 -210
rect 122 -209 126 -196
rect 138 -200 142 -197
rect 129 -204 133 -200
rect 137 -204 142 -200
rect 129 -205 142 -204
rect 122 -213 136 -209
rect 140 -213 141 -209
rect -127 -219 -124 -218
rect -129 -222 -124 -219
rect -120 -222 -114 -218
rect -110 -222 -46 -218
rect -42 -222 7 -218
rect 11 -222 38 -218
rect 42 -222 91 -218
rect 95 -222 108 -218
rect 112 -222 118 -218
rect 122 -222 146 -218
rect -129 -224 146 -222
rect -142 -226 146 -224
rect -142 -227 -125 -226
rect -142 -228 -126 -227
rect -37 -228 7 -226
rect -37 -232 -31 -228
rect -27 -232 -3 -228
rect 1 -232 7 -228
rect -33 -240 -27 -232
rect -33 -244 -32 -240
rect -28 -244 -27 -240
rect -22 -240 -18 -239
rect -13 -240 -7 -232
rect -13 -244 -12 -240
rect -8 -244 -7 -240
rect -2 -240 3 -237
rect 2 -244 3 -240
rect -141 -257 -74 -254
rect -70 -257 -69 -254
rect -329 -279 -324 -278
rect -360 -285 -359 -281
rect -355 -285 -340 -281
rect -337 -283 -329 -281
rect -325 -283 -324 -279
rect -337 -285 -324 -283
rect -342 -291 -341 -288
rect -364 -292 -341 -291
rect -337 -291 -336 -288
rect -337 -292 -330 -291
rect -364 -295 -330 -292
rect -326 -295 -320 -291
rect -364 -296 -320 -295
rect -817 -301 -649 -298
rect -817 -302 -689 -301
rect -511 -302 -496 -298
rect -692 -305 -689 -302
rect -488 -299 -320 -296
rect -161 -293 -156 -273
rect -64 -285 -60 -245
rect -22 -247 -18 -244
rect -2 -245 3 -244
rect -22 -251 -5 -247
rect -52 -279 -49 -252
rect -33 -263 -29 -253
rect -25 -258 -20 -254
rect -9 -255 -5 -251
rect -25 -266 -19 -262
rect -15 -266 -12 -262
rect -25 -272 -21 -266
rect -9 -270 -5 -259
rect -38 -275 -21 -272
rect -17 -274 -5 -270
rect -1 -249 3 -245
rect -1 -252 11 -249
rect -17 -278 -13 -274
rect -1 -275 3 -252
rect 19 -273 22 -258
rect -2 -276 3 -275
rect -33 -282 -32 -278
rect -28 -282 -13 -278
rect -10 -280 -2 -278
rect 2 -280 3 -276
rect -10 -282 3 -280
rect -15 -288 -14 -285
rect -64 -290 -60 -289
rect -37 -289 -14 -288
rect -10 -288 -9 -285
rect 18 -286 23 -273
rect -10 -289 -3 -288
rect -37 -292 -3 -289
rect 1 -292 7 -288
rect -37 -293 7 -292
rect -161 -296 7 -293
rect -161 -297 -37 -296
rect -488 -300 -362 -299
rect -32 -300 -29 -296
rect -365 -303 -362 -300
rect -817 -309 -511 -305
rect -817 -313 -781 -309
rect -777 -313 -767 -309
rect -763 -313 -753 -309
rect -749 -312 -670 -309
rect -749 -313 -686 -312
rect -817 -424 -813 -313
rect -783 -333 -779 -326
rect -783 -334 -778 -333
rect -783 -338 -782 -334
rect -775 -334 -771 -313
rect -768 -319 -755 -318
rect -768 -323 -765 -319
rect -761 -323 -759 -319
rect -768 -324 -755 -323
rect -768 -331 -762 -324
rect -752 -330 -748 -313
rect -682 -313 -670 -312
rect -666 -312 -586 -309
rect -666 -313 -602 -312
rect -705 -324 -693 -318
rect -686 -319 -682 -316
rect -598 -313 -586 -312
rect -582 -313 -549 -309
rect -545 -313 -535 -309
rect -531 -313 -521 -309
rect -517 -313 -511 -309
rect -488 -307 -182 -303
rect -488 -311 -452 -307
rect -448 -311 -438 -307
rect -434 -311 -424 -307
rect -420 -310 -341 -307
rect -420 -311 -357 -310
rect -672 -322 -650 -318
rect -646 -322 -645 -318
rect -621 -319 -609 -318
rect -633 -322 -616 -319
rect -672 -323 -668 -322
rect -686 -324 -682 -323
rect -705 -327 -700 -324
rect -705 -328 -704 -327
rect -775 -338 -772 -334
rect -768 -338 -767 -334
rect -763 -338 -762 -334
rect -758 -338 -757 -334
rect -752 -335 -748 -334
rect -713 -331 -704 -328
rect -679 -327 -668 -323
rect -679 -331 -675 -327
rect -661 -330 -660 -326
rect -656 -330 -645 -326
rect -783 -339 -778 -338
rect -783 -347 -779 -339
rect -763 -343 -757 -338
rect -776 -347 -775 -343
rect -771 -347 -757 -343
rect -751 -345 -747 -342
rect -713 -345 -710 -331
rect -705 -332 -700 -331
rect -696 -333 -675 -331
rect -783 -356 -779 -351
rect -783 -357 -778 -356
rect -783 -361 -782 -357
rect -778 -361 -771 -358
rect -783 -364 -771 -361
rect -767 -360 -763 -347
rect -704 -337 -696 -336
rect -692 -335 -675 -333
rect -704 -340 -692 -337
rect -751 -351 -747 -349
rect -760 -355 -756 -351
rect -752 -355 -747 -351
rect -760 -356 -747 -355
rect -704 -352 -700 -340
rect -679 -342 -675 -335
rect -671 -337 -670 -333
rect -666 -334 -665 -333
rect -666 -337 -654 -334
rect -671 -338 -654 -337
rect -658 -341 -654 -338
rect -658 -342 -653 -341
rect -690 -348 -684 -343
rect -679 -346 -667 -342
rect -663 -346 -662 -342
rect -658 -346 -657 -342
rect -690 -350 -688 -348
rect -697 -352 -688 -350
rect -658 -347 -653 -346
rect -649 -346 -645 -330
rect -658 -351 -654 -347
rect -697 -356 -684 -352
rect -678 -355 -654 -351
rect -649 -350 -647 -346
rect -704 -357 -700 -356
rect -678 -357 -674 -355
rect -767 -364 -753 -360
rect -749 -364 -748 -360
rect -691 -364 -690 -360
rect -686 -364 -685 -360
rect -649 -359 -645 -350
rect -678 -362 -674 -361
rect -669 -363 -668 -359
rect -664 -363 -645 -359
rect -633 -362 -630 -322
rect -621 -323 -616 -322
rect -612 -323 -609 -319
rect -621 -324 -609 -323
rect -602 -319 -598 -316
rect -588 -322 -566 -318
rect -562 -322 -561 -318
rect -588 -323 -584 -322
rect -602 -324 -598 -323
rect -621 -327 -616 -324
rect -621 -331 -620 -327
rect -595 -327 -584 -323
rect -595 -331 -591 -327
rect -577 -330 -576 -326
rect -572 -330 -561 -326
rect -621 -332 -616 -331
rect -612 -333 -591 -331
rect -620 -337 -612 -336
rect -608 -335 -591 -333
rect -620 -340 -608 -337
rect -620 -352 -616 -340
rect -595 -342 -591 -335
rect -587 -337 -586 -333
rect -582 -334 -581 -333
rect -582 -337 -570 -334
rect -587 -338 -570 -337
rect -574 -341 -570 -338
rect -574 -342 -569 -341
rect -606 -348 -600 -343
rect -595 -346 -583 -342
rect -579 -346 -578 -342
rect -574 -346 -573 -342
rect -606 -350 -604 -348
rect -613 -352 -604 -350
rect -574 -347 -569 -346
rect -574 -351 -570 -347
rect -613 -356 -600 -352
rect -594 -355 -570 -351
rect -620 -357 -616 -356
rect -594 -357 -590 -355
rect -691 -369 -685 -364
rect -607 -364 -606 -360
rect -602 -364 -601 -360
rect -565 -359 -561 -330
rect -551 -333 -547 -326
rect -551 -334 -546 -333
rect -551 -338 -550 -334
rect -543 -334 -539 -313
rect -536 -319 -523 -318
rect -536 -323 -533 -319
rect -529 -323 -527 -319
rect -536 -324 -523 -323
rect -536 -331 -530 -324
rect -520 -330 -516 -313
rect -543 -338 -540 -334
rect -536 -338 -535 -334
rect -531 -338 -530 -334
rect -526 -338 -525 -334
rect -520 -335 -516 -334
rect -551 -339 -546 -338
rect -551 -347 -547 -339
rect -531 -343 -525 -338
rect -544 -347 -543 -343
rect -539 -347 -525 -343
rect -519 -344 -515 -342
rect -594 -362 -590 -361
rect -585 -363 -584 -359
rect -580 -363 -561 -359
rect -557 -350 -547 -347
rect -557 -362 -554 -350
rect -607 -369 -601 -364
rect -551 -356 -547 -350
rect -551 -357 -546 -356
rect -551 -361 -550 -357
rect -546 -361 -539 -358
rect -551 -364 -539 -361
rect -535 -360 -531 -347
rect -519 -351 -515 -348
rect -528 -355 -524 -351
rect -520 -355 -515 -351
rect -528 -356 -515 -355
rect -535 -364 -521 -360
rect -517 -364 -516 -360
rect -784 -373 -781 -369
rect -777 -373 -771 -369
rect -767 -373 -703 -369
rect -699 -373 -650 -369
rect -646 -373 -619 -369
rect -615 -373 -566 -369
rect -562 -373 -549 -369
rect -545 -373 -539 -369
rect -535 -373 -516 -369
rect -784 -376 -516 -373
rect -784 -377 -511 -376
rect -694 -379 -650 -377
rect -694 -383 -688 -379
rect -684 -383 -660 -379
rect -656 -383 -650 -379
rect -690 -391 -684 -383
rect -690 -395 -689 -391
rect -685 -395 -684 -391
rect -679 -391 -675 -390
rect -670 -391 -664 -383
rect -563 -386 -522 -383
rect -670 -395 -669 -391
rect -665 -395 -664 -391
rect -659 -391 -654 -388
rect -655 -395 -654 -391
rect -679 -398 -675 -395
rect -659 -396 -654 -395
rect -679 -402 -662 -398
rect -690 -414 -686 -404
rect -682 -409 -677 -405
rect -666 -406 -662 -402
rect -682 -417 -676 -413
rect -672 -417 -669 -413
rect -818 -444 -813 -424
rect -682 -423 -678 -417
rect -666 -421 -662 -410
rect -695 -426 -678 -423
rect -674 -425 -662 -421
rect -674 -429 -670 -425
rect -658 -426 -654 -396
rect -566 -404 -543 -401
rect -538 -404 -537 -401
rect -659 -427 -654 -426
rect -690 -433 -689 -429
rect -685 -433 -670 -429
rect -667 -431 -659 -429
rect -655 -431 -654 -427
rect -667 -433 -654 -431
rect -672 -439 -671 -436
rect -694 -440 -671 -439
rect -667 -439 -666 -436
rect -667 -440 -660 -439
rect -694 -443 -660 -440
rect -656 -443 -650 -439
rect -694 -444 -650 -443
rect -818 -447 -650 -444
rect -818 -448 -694 -447
rect -525 -487 -522 -386
rect -513 -405 -497 -401
rect -488 -422 -484 -311
rect -454 -331 -450 -324
rect -454 -332 -449 -331
rect -454 -336 -453 -332
rect -446 -332 -442 -311
rect -439 -317 -426 -316
rect -439 -321 -436 -317
rect -432 -321 -430 -317
rect -439 -322 -426 -321
rect -439 -329 -433 -322
rect -423 -328 -419 -311
rect -353 -311 -341 -310
rect -337 -310 -257 -307
rect -337 -311 -273 -310
rect -376 -322 -364 -316
rect -357 -317 -353 -314
rect -269 -311 -257 -310
rect -253 -311 -220 -307
rect -216 -311 -206 -307
rect -202 -311 -192 -307
rect -188 -311 -182 -307
rect -161 -304 145 -300
rect -161 -308 -125 -304
rect -121 -308 -111 -304
rect -107 -308 -97 -304
rect -93 -307 -14 -304
rect -93 -308 -30 -307
rect -343 -320 -321 -316
rect -317 -320 -316 -316
rect -292 -317 -280 -316
rect -343 -321 -339 -320
rect -357 -322 -353 -321
rect -376 -325 -371 -322
rect -376 -326 -375 -325
rect -446 -336 -443 -332
rect -439 -336 -438 -332
rect -434 -336 -433 -332
rect -429 -336 -428 -332
rect -423 -333 -419 -332
rect -384 -329 -375 -326
rect -350 -325 -339 -321
rect -292 -321 -287 -317
rect -283 -321 -280 -317
rect -292 -322 -280 -321
rect -273 -317 -269 -314
rect -259 -320 -237 -316
rect -233 -320 -232 -316
rect -259 -321 -255 -320
rect -273 -322 -269 -321
rect -350 -329 -346 -325
rect -332 -328 -331 -324
rect -327 -328 -316 -324
rect -454 -337 -449 -336
rect -454 -345 -450 -337
rect -434 -341 -428 -336
rect -447 -345 -446 -341
rect -442 -345 -428 -341
rect -422 -343 -418 -340
rect -454 -354 -450 -349
rect -454 -355 -449 -354
rect -454 -359 -453 -355
rect -449 -359 -442 -356
rect -454 -362 -442 -359
rect -438 -358 -434 -345
rect -422 -349 -418 -347
rect -431 -353 -427 -349
rect -423 -353 -418 -349
rect -431 -354 -418 -353
rect -438 -362 -424 -358
rect -420 -362 -419 -358
rect -394 -360 -391 -340
rect -384 -343 -381 -329
rect -376 -330 -371 -329
rect -367 -331 -346 -329
rect -375 -335 -367 -334
rect -363 -333 -346 -331
rect -375 -338 -363 -335
rect -375 -350 -371 -338
rect -350 -340 -346 -333
rect -342 -335 -341 -331
rect -337 -332 -336 -331
rect -337 -335 -325 -332
rect -342 -336 -325 -335
rect -329 -339 -325 -336
rect -329 -340 -324 -339
rect -361 -346 -355 -341
rect -350 -344 -338 -340
rect -334 -344 -333 -340
rect -329 -344 -328 -340
rect -361 -348 -359 -346
rect -368 -350 -359 -348
rect -329 -345 -324 -344
rect -320 -344 -316 -328
rect -292 -325 -287 -322
rect -292 -329 -291 -325
rect -266 -325 -255 -321
rect -266 -329 -262 -325
rect -248 -328 -247 -324
rect -243 -328 -232 -324
rect -292 -330 -287 -329
rect -283 -331 -262 -329
rect -291 -335 -283 -334
rect -279 -333 -262 -331
rect -291 -338 -279 -335
rect -329 -349 -325 -345
rect -368 -354 -355 -350
rect -349 -353 -325 -349
rect -320 -348 -318 -344
rect -375 -355 -371 -354
rect -349 -355 -345 -353
rect -362 -362 -361 -358
rect -357 -362 -356 -358
rect -320 -357 -316 -348
rect -291 -350 -287 -338
rect -266 -340 -262 -333
rect -258 -335 -257 -331
rect -253 -332 -252 -331
rect -253 -335 -241 -332
rect -258 -336 -241 -335
rect -245 -339 -241 -336
rect -245 -340 -240 -339
rect -277 -346 -271 -341
rect -266 -344 -254 -340
rect -250 -344 -249 -340
rect -245 -344 -244 -340
rect -277 -348 -275 -346
rect -284 -350 -275 -348
rect -245 -345 -240 -344
rect -245 -349 -241 -345
rect -284 -354 -271 -350
rect -265 -353 -241 -349
rect -291 -355 -287 -354
rect -265 -355 -261 -353
rect -349 -360 -345 -359
rect -340 -361 -339 -357
rect -335 -361 -316 -357
rect -362 -367 -356 -362
rect -278 -362 -277 -358
rect -273 -362 -272 -358
rect -236 -357 -232 -328
rect -222 -331 -218 -324
rect -222 -332 -217 -331
rect -222 -336 -221 -332
rect -214 -332 -210 -311
rect -207 -317 -194 -316
rect -207 -321 -204 -317
rect -200 -321 -198 -317
rect -207 -322 -194 -321
rect -207 -329 -201 -322
rect -191 -328 -187 -311
rect -214 -336 -211 -332
rect -207 -336 -206 -332
rect -202 -336 -201 -332
rect -197 -336 -196 -332
rect -191 -333 -187 -332
rect -222 -337 -217 -336
rect -222 -345 -218 -337
rect -202 -341 -196 -336
rect -215 -345 -214 -341
rect -210 -345 -196 -341
rect -190 -342 -186 -340
rect -265 -360 -261 -359
rect -256 -361 -255 -357
rect -251 -361 -232 -357
rect -228 -348 -218 -345
rect -228 -360 -225 -348
rect -278 -367 -272 -362
rect -222 -354 -218 -348
rect -222 -355 -217 -354
rect -222 -359 -221 -355
rect -217 -359 -210 -356
rect -222 -362 -210 -359
rect -206 -358 -202 -345
rect -190 -349 -186 -346
rect -199 -353 -195 -349
rect -191 -353 -186 -349
rect -199 -354 -186 -353
rect -206 -362 -192 -358
rect -188 -362 -187 -358
rect -455 -371 -452 -367
rect -448 -371 -442 -367
rect -438 -371 -374 -367
rect -370 -371 -321 -367
rect -317 -371 -290 -367
rect -286 -371 -237 -367
rect -233 -371 -220 -367
rect -216 -371 -210 -367
rect -206 -371 -182 -367
rect -474 -374 -189 -371
rect -455 -375 -189 -374
rect -185 -375 -182 -371
rect -365 -377 -321 -375
rect -365 -381 -359 -377
rect -355 -381 -331 -377
rect -327 -381 -321 -377
rect -394 -386 -391 -384
rect -361 -389 -355 -381
rect -394 -404 -391 -390
rect -361 -393 -360 -389
rect -356 -393 -355 -389
rect -350 -389 -346 -388
rect -341 -389 -335 -381
rect -341 -393 -340 -389
rect -336 -393 -335 -389
rect -330 -389 -325 -386
rect -326 -393 -325 -389
rect -350 -396 -346 -393
rect -330 -394 -325 -393
rect -350 -400 -333 -396
rect -489 -442 -484 -422
rect -422 -408 -394 -405
rect -422 -434 -418 -408
rect -361 -412 -357 -402
rect -353 -407 -348 -403
rect -337 -404 -333 -400
rect -353 -415 -347 -411
rect -343 -415 -340 -411
rect -353 -421 -349 -415
rect -337 -419 -333 -408
rect -366 -424 -349 -421
rect -345 -423 -333 -419
rect -345 -427 -341 -423
rect -329 -424 -325 -394
rect -298 -398 -216 -393
rect -161 -419 -157 -308
rect -127 -328 -123 -321
rect -127 -329 -122 -328
rect -127 -333 -126 -329
rect -119 -329 -115 -308
rect -112 -314 -99 -313
rect -112 -318 -109 -314
rect -105 -318 -103 -314
rect -112 -319 -99 -318
rect -112 -326 -106 -319
rect -96 -325 -92 -308
rect -26 -308 -14 -307
rect -10 -307 70 -304
rect -10 -308 54 -307
rect -49 -319 -37 -313
rect -30 -314 -26 -311
rect 58 -308 70 -307
rect 74 -308 107 -304
rect 111 -308 121 -304
rect 125 -308 135 -304
rect 139 -308 145 -304
rect -16 -317 6 -313
rect 10 -317 11 -313
rect 35 -314 47 -313
rect -16 -318 -12 -317
rect -30 -319 -26 -318
rect -49 -322 -44 -319
rect -49 -323 -48 -322
rect -119 -333 -116 -329
rect -112 -333 -111 -329
rect -107 -333 -106 -329
rect -102 -333 -101 -329
rect -96 -330 -92 -329
rect -57 -326 -48 -323
rect -23 -322 -12 -318
rect 35 -318 40 -314
rect 44 -318 47 -314
rect 35 -319 47 -318
rect 54 -314 58 -311
rect 68 -317 90 -313
rect 94 -317 95 -313
rect 68 -318 72 -317
rect 54 -319 58 -318
rect -23 -326 -19 -322
rect -5 -325 -4 -321
rect 0 -325 11 -321
rect -127 -334 -122 -333
rect -127 -342 -123 -334
rect -107 -338 -101 -333
rect -120 -342 -119 -338
rect -115 -342 -101 -338
rect -95 -340 -91 -337
rect -57 -340 -54 -326
rect -49 -327 -44 -326
rect -40 -328 -19 -326
rect -127 -351 -123 -346
rect -127 -352 -122 -351
rect -127 -356 -126 -352
rect -122 -356 -115 -353
rect -127 -359 -115 -356
rect -111 -355 -107 -342
rect -48 -332 -40 -331
rect -36 -330 -19 -328
rect -48 -335 -36 -332
rect -95 -346 -91 -344
rect -104 -350 -100 -346
rect -96 -350 -91 -346
rect -104 -351 -91 -350
rect -48 -347 -44 -335
rect -23 -337 -19 -330
rect -15 -332 -14 -328
rect -10 -329 -9 -328
rect -10 -332 2 -329
rect -15 -333 2 -332
rect -2 -336 2 -333
rect -2 -337 3 -336
rect -34 -343 -28 -338
rect -23 -341 -11 -337
rect -7 -341 -6 -337
rect -2 -341 -1 -337
rect -34 -345 -32 -343
rect -48 -352 -44 -351
rect -41 -347 -32 -345
rect -2 -342 3 -341
rect 7 -341 11 -325
rect 35 -322 40 -319
rect 35 -326 36 -322
rect 61 -322 72 -318
rect 61 -326 65 -322
rect 79 -325 80 -321
rect 84 -325 95 -321
rect 35 -327 40 -326
rect 44 -328 65 -326
rect 36 -332 44 -331
rect 48 -330 65 -328
rect 36 -335 48 -332
rect -2 -346 2 -342
rect -41 -351 -28 -347
rect -22 -350 2 -346
rect 7 -345 9 -341
rect -111 -359 -97 -355
rect -93 -359 -92 -355
rect -41 -356 -38 -351
rect -22 -352 -18 -350
rect -52 -360 -38 -356
rect -35 -359 -34 -355
rect -30 -359 -29 -355
rect 7 -354 11 -345
rect 36 -347 40 -335
rect 61 -337 65 -330
rect 69 -332 70 -328
rect 74 -329 75 -328
rect 74 -332 86 -329
rect 69 -333 86 -332
rect 82 -336 86 -333
rect 82 -337 87 -336
rect 50 -343 56 -338
rect 61 -341 73 -337
rect 77 -341 78 -337
rect 82 -341 83 -337
rect 50 -345 52 -343
rect 43 -347 52 -345
rect 82 -342 87 -341
rect 82 -346 86 -342
rect 43 -351 56 -347
rect 62 -350 86 -346
rect 36 -352 40 -351
rect 62 -352 66 -350
rect -22 -357 -18 -356
rect -13 -358 -12 -354
rect -8 -358 11 -354
rect -52 -364 -48 -360
rect -35 -364 -29 -359
rect 49 -359 50 -355
rect 54 -359 55 -355
rect 91 -354 95 -325
rect 105 -328 109 -321
rect 105 -329 110 -328
rect 105 -333 106 -329
rect 113 -329 117 -308
rect 120 -314 133 -313
rect 120 -318 123 -314
rect 127 -318 129 -314
rect 120 -319 133 -318
rect 120 -326 126 -319
rect 136 -325 140 -308
rect 113 -333 116 -329
rect 120 -333 121 -329
rect 125 -333 126 -329
rect 130 -333 131 -329
rect 136 -330 140 -329
rect 105 -334 110 -333
rect 105 -342 109 -334
rect 125 -338 131 -333
rect 112 -342 113 -338
rect 117 -342 131 -338
rect 137 -339 141 -337
rect 62 -357 66 -356
rect 71 -358 72 -354
rect 76 -358 95 -354
rect 99 -345 109 -342
rect 99 -357 102 -345
rect 49 -364 55 -359
rect 105 -351 109 -345
rect 105 -352 110 -351
rect 105 -356 106 -352
rect 110 -356 117 -353
rect 105 -359 117 -356
rect 121 -355 125 -342
rect 137 -346 141 -343
rect 128 -350 132 -346
rect 136 -350 141 -346
rect 128 -351 141 -350
rect 121 -359 135 -355
rect 139 -359 140 -355
rect -128 -367 -125 -364
rect -129 -368 -125 -367
rect -121 -368 -115 -364
rect -111 -368 -47 -364
rect -43 -368 6 -364
rect 10 -368 37 -364
rect 41 -368 90 -364
rect 94 -368 107 -364
rect 111 -368 117 -364
rect 121 -368 145 -364
rect -129 -370 145 -368
rect -148 -371 145 -370
rect -145 -372 145 -371
rect -145 -373 -126 -372
rect -38 -374 6 -372
rect -38 -378 -32 -374
rect -28 -378 -4 -374
rect 0 -378 6 -374
rect -91 -380 -87 -379
rect -147 -398 -118 -393
rect -330 -425 -325 -424
rect -361 -431 -360 -427
rect -356 -431 -341 -427
rect -338 -429 -330 -427
rect -326 -427 -325 -425
rect -326 -429 -321 -427
rect -338 -431 -321 -429
rect -343 -437 -342 -434
rect -365 -438 -342 -437
rect -338 -437 -337 -434
rect -338 -438 -331 -437
rect -365 -441 -331 -438
rect -327 -441 -321 -437
rect -365 -442 -321 -441
rect -489 -445 -321 -442
rect -162 -439 -157 -419
rect -91 -421 -87 -384
rect -34 -386 -28 -378
rect -34 -390 -33 -386
rect -29 -390 -28 -386
rect -23 -386 -19 -385
rect -14 -386 -8 -378
rect -14 -390 -13 -386
rect -9 -390 -8 -386
rect -3 -386 2 -383
rect 1 -390 2 -386
rect -23 -393 -19 -390
rect -3 -391 2 -390
rect -23 -397 -6 -393
rect -34 -409 -30 -399
rect -26 -404 -21 -400
rect -10 -401 -6 -397
rect -26 -412 -20 -408
rect -16 -412 -13 -408
rect -26 -418 -22 -412
rect -10 -416 -6 -405
rect -39 -421 -22 -418
rect -18 -420 -6 -416
rect -2 -396 14 -391
rect -18 -424 -14 -420
rect -2 -421 2 -396
rect -3 -422 2 -421
rect -34 -428 -33 -424
rect -29 -428 -14 -424
rect -11 -426 -3 -424
rect 1 -426 2 -422
rect -11 -428 2 -426
rect -16 -434 -15 -431
rect -38 -435 -15 -434
rect -11 -434 -10 -431
rect -11 -435 -4 -434
rect -38 -438 -4 -435
rect 0 -438 6 -434
rect -38 -439 6 -438
rect -162 -442 6 -439
rect -162 -443 -38 -442
rect -489 -446 -365 -445
rect -376 -453 -372 -446
rect -493 -455 -449 -453
rect -400 -455 -356 -453
rect -313 -455 -269 -453
rect -493 -457 -269 -455
rect -493 -461 -487 -457
rect -483 -458 -394 -457
rect -483 -461 -449 -458
rect -400 -461 -394 -458
rect -390 -458 -307 -457
rect -390 -461 -356 -458
rect -313 -461 -307 -458
rect -303 -461 -269 -457
rect -479 -469 -473 -461
rect -479 -473 -478 -469
rect -474 -473 -473 -469
rect -468 -467 -464 -466
rect -459 -467 -453 -461
rect -418 -467 -407 -464
rect -459 -471 -458 -467
rect -454 -471 -453 -467
rect -489 -474 -484 -473
rect -489 -478 -488 -474
rect -468 -474 -464 -471
rect -489 -481 -484 -478
rect -489 -485 -488 -481
rect -489 -486 -484 -485
rect -481 -478 -468 -476
rect -481 -480 -464 -478
rect -457 -478 -426 -474
rect -489 -487 -485 -486
rect -525 -491 -485 -487
rect -489 -504 -485 -491
rect -481 -491 -477 -480
rect -466 -487 -461 -483
rect -457 -487 -453 -478
rect -474 -495 -471 -491
rect -467 -495 -460 -491
rect -481 -499 -477 -495
rect -481 -503 -469 -499
rect -465 -500 -460 -495
rect -489 -505 -484 -504
rect -489 -509 -488 -505
rect -484 -509 -477 -506
rect -489 -512 -477 -509
rect -473 -507 -469 -503
rect -466 -504 -450 -500
rect -473 -511 -458 -507
rect -454 -511 -453 -507
rect -430 -511 -426 -478
rect -410 -477 -407 -467
rect -386 -469 -380 -461
rect -386 -473 -385 -469
rect -381 -473 -380 -469
rect -375 -467 -371 -466
rect -366 -467 -360 -461
rect -366 -471 -365 -467
rect -361 -471 -360 -467
rect -299 -469 -293 -461
rect -320 -470 -304 -469
rect -396 -474 -391 -473
rect -396 -477 -395 -474
rect -410 -478 -395 -477
rect -375 -474 -371 -471
rect -410 -480 -391 -478
rect -396 -481 -391 -480
rect -396 -485 -395 -481
rect -396 -486 -391 -485
rect -388 -478 -375 -476
rect -388 -480 -371 -478
rect -396 -504 -392 -486
rect -388 -491 -384 -480
rect -364 -483 -360 -474
rect -316 -474 -304 -470
rect -299 -473 -298 -469
rect -294 -473 -293 -469
rect -288 -467 -284 -466
rect -279 -467 -273 -461
rect -279 -471 -278 -467
rect -274 -471 -273 -467
rect -316 -475 -308 -474
rect -309 -478 -308 -475
rect -288 -474 -284 -471
rect -309 -481 -304 -478
rect -373 -487 -368 -483
rect -364 -487 -353 -483
rect -309 -485 -308 -481
rect -309 -486 -304 -485
rect -301 -478 -288 -476
rect -301 -480 -284 -478
rect -381 -495 -378 -491
rect -374 -495 -367 -491
rect -388 -499 -384 -495
rect -388 -503 -376 -499
rect -396 -505 -391 -504
rect -396 -509 -395 -505
rect -391 -509 -384 -506
rect -396 -512 -384 -509
rect -380 -507 -376 -503
rect -372 -500 -367 -495
rect -372 -504 -357 -500
rect -309 -504 -305 -486
rect -301 -491 -297 -480
rect -277 -483 -273 -474
rect -286 -487 -281 -483
rect -277 -487 -264 -483
rect -294 -495 -291 -491
rect -287 -495 -280 -491
rect -301 -499 -297 -495
rect -301 -503 -289 -499
rect -309 -505 -304 -504
rect -380 -511 -365 -507
rect -361 -511 -360 -507
rect -309 -509 -308 -505
rect -304 -509 -297 -506
rect -309 -512 -297 -509
rect -293 -507 -289 -503
rect -285 -501 -280 -495
rect -285 -504 -272 -501
rect -293 -511 -278 -507
rect -274 -511 -273 -507
rect -493 -521 -487 -517
rect -483 -521 -477 -517
rect -473 -521 -449 -517
rect -400 -521 -394 -517
rect -390 -521 -384 -517
rect -380 -521 -356 -517
rect -499 -522 -356 -521
rect -313 -521 -307 -517
rect -303 -521 -297 -517
rect -293 -521 -269 -517
rect -313 -522 -269 -521
rect -499 -524 -269 -522
rect -493 -525 -449 -524
rect -400 -525 -269 -524
<< metal2 >>
rect -30 -39 50 -36
rect -30 -45 -27 -39
rect -69 -48 -27 -45
rect 46 -46 49 -39
rect 70 -41 129 -38
rect 3 -49 24 -46
rect 50 -49 76 -46
rect 80 -49 81 -46
rect 126 -47 129 -41
rect 150 -46 169 -43
rect 126 -50 133 -47
rect 150 -51 153 -46
rect 173 -45 212 -44
rect 173 -47 208 -45
rect -54 -59 -42 -56
rect -737 -81 -708 -77
rect -801 -85 -734 -81
rect -801 -227 -796 -85
rect -727 -92 -474 -88
rect -786 -150 -782 -99
rect -727 -127 -722 -92
rect -479 -96 -475 -92
rect -709 -105 -708 -102
rect -704 -105 -620 -102
rect -616 -105 -527 -102
rect -344 -106 -340 -72
rect -302 -91 -54 -87
rect -302 -95 -298 -91
rect -245 -103 -156 -100
rect -247 -104 -156 -103
rect -152 -104 -69 -100
rect -623 -123 -479 -120
rect -297 -121 -150 -118
rect -728 -131 -716 -127
rect -623 -127 -620 -123
rect -153 -125 -150 -121
rect -711 -131 -700 -127
rect -571 -132 -570 -129
rect -787 -152 -782 -150
rect -787 -188 -783 -152
rect -643 -153 -595 -150
rect -643 -154 -586 -153
rect -598 -157 -586 -154
rect -573 -163 -570 -132
rect -530 -137 -527 -131
rect -249 -129 -245 -126
rect -530 -140 -479 -137
rect -249 -137 -246 -129
rect -297 -140 -246 -137
rect -153 -129 -152 -125
rect -135 -127 -116 -123
rect -58 -125 -54 -91
rect -45 -98 -42 -59
rect 18 -59 100 -56
rect 163 -56 222 -53
rect 133 -61 136 -58
rect 133 -64 191 -61
rect 122 -83 126 -65
rect 3 -87 126 -83
rect 2 -91 6 -87
rect 122 -88 126 -87
rect 2 -109 5 -91
rect 12 -94 29 -91
rect 10 -96 15 -94
rect 14 -97 15 -96
rect 26 -97 29 -94
rect 26 -100 74 -97
rect 137 -102 195 -99
rect 22 -107 104 -104
rect 137 -105 140 -102
rect 1 -113 7 -109
rect 167 -110 226 -107
rect 1 -116 3 -113
rect 7 -117 28 -114
rect 54 -117 80 -114
rect 84 -117 96 -114
rect 129 -116 137 -113
rect 50 -123 53 -117
rect 129 -121 132 -116
rect 177 -118 212 -116
rect 177 -119 216 -118
rect 76 -124 132 -121
rect -72 -129 -64 -125
rect -59 -127 -54 -125
rect -59 -129 68 -127
rect 137 -128 168 -127
rect -252 -148 -249 -140
rect -325 -151 -314 -149
rect -252 -151 -238 -148
rect -325 -152 -320 -151
rect -544 -155 -320 -152
rect -316 -155 -314 -151
rect -544 -156 -314 -155
rect -214 -157 -211 -130
rect -152 -139 -149 -129
rect -58 -130 68 -129
rect 81 -130 168 -128
rect -45 -131 168 -130
rect 62 -134 86 -131
rect 154 -139 158 -138
rect -152 -143 158 -139
rect -199 -151 -140 -148
rect -309 -160 -211 -157
rect -112 -151 150 -148
rect -126 -155 -122 -152
rect -126 -158 -59 -155
rect -621 -164 -568 -163
rect -703 -167 -568 -164
rect -309 -165 -305 -160
rect -703 -173 -700 -167
rect -754 -176 -689 -173
rect -787 -192 -746 -188
rect -750 -199 -746 -192
rect -797 -231 -796 -227
rect -789 -201 -786 -200
rect -789 -204 -782 -201
rect -789 -269 -786 -204
rect -746 -203 -713 -200
rect -693 -200 -690 -176
rect -611 -176 -526 -173
rect -522 -176 -501 -173
rect -425 -174 -360 -171
rect -642 -204 -609 -201
rect -629 -208 -626 -204
rect -517 -208 -514 -202
rect -629 -211 -514 -208
rect -553 -220 -552 -217
rect -555 -268 -552 -220
rect -504 -226 -501 -176
rect -364 -177 -360 -174
rect -309 -177 -306 -165
rect -63 -168 -59 -158
rect -302 -171 -282 -169
rect -302 -172 -286 -171
rect -302 -176 -301 -172
rect -297 -175 -286 -172
rect -282 -174 -197 -171
rect -98 -171 -33 -168
rect -297 -176 -282 -175
rect -302 -177 -294 -176
rect -364 -180 -306 -177
rect -460 -202 -453 -199
rect -510 -230 -476 -226
rect -516 -231 -476 -230
rect -789 -272 -695 -269
rect -685 -271 -542 -268
rect -698 -276 -695 -272
rect -547 -302 -516 -298
rect -566 -303 -542 -302
rect -609 -306 -542 -303
rect -609 -307 -606 -306
rect -665 -310 -606 -307
rect -665 -319 -661 -310
rect -755 -322 -661 -319
rect -790 -350 -783 -347
rect -790 -415 -787 -350
rect -747 -349 -714 -346
rect -694 -346 -691 -322
rect -612 -322 -527 -319
rect -733 -384 -730 -349
rect -643 -350 -610 -347
rect -630 -354 -627 -350
rect -518 -354 -515 -348
rect -630 -357 -515 -354
rect -554 -366 -553 -363
rect -633 -382 -630 -366
rect -733 -388 -640 -384
rect -634 -385 -567 -382
rect -645 -401 -640 -388
rect -645 -405 -572 -401
rect -556 -414 -553 -366
rect -503 -370 -500 -231
rect -492 -254 -471 -250
rect -460 -267 -457 -202
rect -417 -201 -384 -198
rect -364 -198 -361 -180
rect -225 -182 -67 -179
rect -399 -250 -395 -201
rect -313 -202 -280 -199
rect -300 -206 -297 -202
rect -188 -206 -185 -200
rect -300 -209 -185 -206
rect -133 -199 -126 -196
rect -224 -218 -223 -215
rect -226 -266 -223 -218
rect -183 -228 -149 -224
rect -189 -229 -149 -228
rect -173 -257 -145 -254
rect -133 -264 -130 -199
rect -90 -198 -57 -195
rect -37 -195 -34 -171
rect 45 -171 130 -168
rect 22 -179 96 -177
rect 22 -180 100 -179
rect -74 -253 -70 -198
rect 14 -199 47 -196
rect 27 -203 30 -199
rect 139 -203 142 -197
rect 27 -206 142 -203
rect -65 -240 -62 -215
rect 103 -215 104 -212
rect -48 -252 11 -249
rect 19 -253 23 -215
rect 101 -263 104 -215
rect -460 -270 -366 -267
rect -356 -269 -213 -266
rect -133 -267 -39 -264
rect -29 -266 114 -263
rect -369 -274 -366 -270
rect -42 -271 -39 -267
rect -71 -278 -51 -275
rect -71 -280 -68 -278
rect -311 -283 -68 -280
rect -54 -279 -51 -278
rect 9 -278 57 -275
rect -54 -283 -52 -279
rect -48 -283 -47 -280
rect -311 -299 -308 -283
rect 9 -287 12 -278
rect -60 -289 12 -287
rect -64 -290 12 -289
rect 18 -296 23 -293
rect -491 -302 -308 -299
rect -282 -300 23 -296
rect -282 -301 -159 -300
rect -281 -317 -276 -301
rect 51 -314 54 -278
rect -426 -320 -361 -317
rect -394 -336 -391 -320
rect -461 -348 -454 -345
rect -508 -371 -478 -370
rect -508 -376 -479 -371
rect -538 -405 -518 -401
rect -790 -418 -696 -415
rect -686 -417 -543 -414
rect -699 -422 -696 -418
rect -507 -519 -501 -376
rect -480 -401 -476 -400
rect -492 -405 -476 -401
rect -480 -426 -476 -405
rect -461 -413 -458 -348
rect -418 -347 -385 -344
rect -365 -344 -362 -320
rect -283 -320 -198 -317
rect -99 -317 -34 -314
rect -403 -394 -400 -347
rect -314 -348 -281 -345
rect -301 -352 -298 -348
rect -189 -352 -186 -346
rect -301 -355 -186 -352
rect -134 -345 -127 -342
rect -394 -360 -391 -359
rect -225 -364 -224 -361
rect -394 -386 -391 -364
rect -403 -398 -304 -394
rect -227 -412 -224 -364
rect -185 -374 -149 -371
rect -211 -398 -152 -393
rect -134 -410 -131 -345
rect -91 -344 -58 -341
rect -38 -341 -35 -317
rect 44 -317 129 -314
rect -71 -380 -67 -344
rect 13 -345 46 -342
rect 26 -349 29 -345
rect 138 -349 141 -343
rect 26 -352 141 -349
rect 102 -361 103 -358
rect -87 -384 -67 -380
rect -71 -385 -67 -384
rect -113 -396 14 -393
rect 20 -396 21 -393
rect -113 -397 21 -396
rect 100 -409 103 -361
rect -461 -416 -367 -413
rect -357 -415 -214 -412
rect -134 -413 -40 -410
rect -30 -412 113 -409
rect -370 -420 -367 -416
rect -43 -417 -40 -413
rect -91 -421 -87 -420
rect -480 -430 -403 -426
rect -406 -434 -403 -430
rect -323 -431 -321 -426
rect -323 -434 -318 -431
rect -422 -463 -418 -438
rect -406 -438 -318 -434
rect -406 -439 -403 -438
rect -91 -470 -87 -425
rect 147 -431 150 -151
rect -316 -473 -87 -470
rect -316 -474 -91 -473
rect 146 -483 150 -431
rect -349 -487 -315 -483
rect -260 -486 150 -483
rect 146 -487 150 -486
rect -319 -491 -315 -487
rect -319 -494 -250 -491
rect -253 -498 -250 -494
rect 154 -498 158 -143
rect -445 -504 -357 -500
rect -352 -504 -272 -501
rect -253 -502 158 -498
rect 165 -512 168 -131
rect -426 -515 168 -512
rect -507 -526 -506 -519
<< metal3 >>
rect -321 -151 -296 -149
rect -321 -155 -320 -151
rect -316 -155 -296 -151
rect -321 -156 -315 -155
rect -302 -170 -296 -155
rect -302 -172 -295 -170
rect -302 -176 -301 -172
rect -297 -176 -295 -172
rect -302 -177 -295 -176
<< ntransistor >>
rect -78 -71 -76 -68
rect -6 -72 -4 -69
rect 33 -72 35 -66
rect 54 -72 56 -66
rect 87 -72 89 -66
rect 108 -72 110 -66
rect 143 -72 145 -66
rect 164 -72 166 -66
rect 197 -72 199 -66
rect 218 -72 220 -66
rect -697 -104 -695 -93
rect -690 -104 -688 -93
rect -677 -104 -675 -95
rect -610 -104 -608 -93
rect -603 -104 -601 -93
rect -590 -104 -588 -95
rect -517 -104 -515 -93
rect -510 -104 -508 -93
rect -497 -104 -495 -95
rect -277 -102 -275 -93
rect -264 -102 -262 -91
rect -257 -102 -255 -91
rect -184 -102 -182 -93
rect -171 -102 -169 -91
rect -164 -102 -162 -91
rect -97 -102 -95 -93
rect -84 -102 -82 -91
rect -77 -102 -75 -91
rect -2 -94 0 -91
rect 37 -97 39 -91
rect 58 -97 60 -91
rect 91 -97 93 -91
rect 112 -97 114 -91
rect 147 -97 149 -91
rect 168 -97 170 -91
rect 201 -97 203 -91
rect 222 -97 224 -91
rect -775 -216 -773 -210
rect -763 -222 -761 -213
rect -756 -222 -754 -213
rect -697 -214 -695 -205
rect -681 -219 -679 -210
rect -671 -219 -669 -210
rect -661 -222 -659 -210
rect -654 -222 -652 -210
rect -613 -214 -611 -205
rect -597 -219 -595 -210
rect -587 -219 -585 -210
rect -577 -222 -575 -210
rect -570 -222 -568 -210
rect -543 -216 -541 -210
rect -531 -222 -529 -213
rect -524 -222 -522 -213
rect -446 -214 -444 -208
rect -434 -220 -432 -211
rect -427 -220 -425 -211
rect -368 -212 -366 -203
rect -352 -217 -350 -208
rect -342 -217 -340 -208
rect -332 -220 -330 -208
rect -325 -220 -323 -208
rect -284 -212 -282 -203
rect -268 -217 -266 -208
rect -258 -217 -256 -208
rect -248 -220 -246 -208
rect -241 -220 -239 -208
rect -214 -214 -212 -208
rect -119 -211 -117 -205
rect -202 -220 -200 -211
rect -195 -220 -193 -211
rect -107 -217 -105 -208
rect -100 -217 -98 -208
rect -41 -209 -39 -200
rect -25 -214 -23 -205
rect -15 -214 -13 -205
rect -5 -217 -3 -205
rect 2 -217 4 -205
rect 43 -209 45 -200
rect 59 -214 61 -205
rect 69 -214 71 -205
rect 79 -217 81 -205
rect 86 -217 88 -205
rect 113 -211 115 -205
rect 125 -217 127 -208
rect 132 -217 134 -208
rect -682 -250 -680 -244
rect -672 -250 -670 -244
rect -662 -250 -660 -244
rect -353 -248 -351 -242
rect -343 -248 -341 -242
rect -333 -248 -331 -242
rect -26 -245 -24 -239
rect -16 -245 -14 -239
rect -6 -245 -4 -239
rect -776 -362 -774 -356
rect -764 -368 -762 -359
rect -757 -368 -755 -359
rect -698 -360 -696 -351
rect -682 -365 -680 -356
rect -672 -365 -670 -356
rect -662 -368 -660 -356
rect -655 -368 -653 -356
rect -614 -360 -612 -351
rect -598 -365 -596 -356
rect -588 -365 -586 -356
rect -578 -368 -576 -356
rect -571 -368 -569 -356
rect -544 -362 -542 -356
rect -532 -368 -530 -359
rect -525 -368 -523 -359
rect -447 -360 -445 -354
rect -435 -366 -433 -357
rect -428 -366 -426 -357
rect -369 -358 -367 -349
rect -353 -363 -351 -354
rect -343 -363 -341 -354
rect -333 -366 -331 -354
rect -326 -366 -324 -354
rect -285 -358 -283 -349
rect -269 -363 -267 -354
rect -259 -363 -257 -354
rect -249 -366 -247 -354
rect -242 -366 -240 -354
rect -215 -360 -213 -354
rect -120 -357 -118 -351
rect -203 -366 -201 -357
rect -196 -366 -194 -357
rect -108 -363 -106 -354
rect -101 -363 -99 -354
rect -42 -355 -40 -346
rect -26 -360 -24 -351
rect -16 -360 -14 -351
rect -6 -363 -4 -351
rect 1 -363 3 -351
rect 42 -355 44 -346
rect 58 -360 60 -351
rect 68 -360 70 -351
rect 78 -363 80 -351
rect 85 -363 87 -351
rect 112 -357 114 -351
rect 124 -363 126 -354
rect 131 -363 133 -354
rect -683 -396 -681 -390
rect -673 -396 -671 -390
rect -663 -396 -661 -390
rect -354 -394 -352 -388
rect -344 -394 -342 -388
rect -334 -394 -332 -388
rect -27 -391 -25 -385
rect -17 -391 -15 -385
rect -7 -391 -5 -385
rect -482 -510 -480 -501
rect -469 -512 -467 -501
rect -462 -512 -460 -501
rect -389 -510 -387 -501
rect -376 -512 -374 -501
rect -369 -512 -367 -501
rect -302 -510 -300 -501
rect -289 -512 -287 -501
rect -282 -512 -280 -501
<< ptransistor >>
rect -78 -35 -76 -29
rect -6 -35 -4 -29
rect 33 -35 35 -29
rect 54 -35 56 -29
rect 87 -35 89 -29
rect 108 -35 110 -29
rect 143 -35 145 -29
rect 164 -35 166 -29
rect 197 -35 199 -29
rect 218 -35 220 -29
rect -697 -139 -695 -126
rect -687 -139 -685 -126
rect -677 -137 -675 -119
rect -610 -139 -608 -126
rect -600 -139 -598 -126
rect -590 -137 -588 -119
rect -517 -139 -515 -126
rect -507 -139 -505 -126
rect -497 -137 -495 -119
rect -277 -135 -275 -117
rect -267 -137 -265 -124
rect -257 -137 -255 -124
rect -184 -135 -182 -117
rect -174 -137 -172 -124
rect -164 -137 -162 -124
rect -97 -135 -95 -117
rect -87 -137 -85 -124
rect -77 -137 -75 -124
rect -2 -134 0 -128
rect 37 -134 39 -128
rect 58 -134 60 -128
rect 91 -134 93 -128
rect 112 -134 114 -128
rect 147 -134 149 -128
rect 168 -134 170 -128
rect 201 -134 203 -128
rect 222 -134 224 -128
rect -775 -193 -773 -181
rect -765 -193 -763 -183
rect -755 -193 -753 -183
rect -689 -192 -687 -165
rect -673 -192 -671 -174
rect -663 -192 -661 -174
rect -653 -192 -651 -165
rect -605 -192 -603 -165
rect -589 -192 -587 -174
rect -579 -192 -577 -174
rect -569 -192 -567 -165
rect -543 -193 -541 -181
rect -533 -193 -531 -183
rect -523 -193 -521 -183
rect -446 -191 -444 -179
rect -436 -191 -434 -181
rect -426 -191 -424 -181
rect -360 -190 -358 -163
rect -344 -190 -342 -172
rect -334 -190 -332 -172
rect -324 -190 -322 -163
rect -276 -190 -274 -163
rect -260 -190 -258 -172
rect -250 -190 -248 -172
rect -240 -190 -238 -163
rect -214 -191 -212 -179
rect -204 -191 -202 -181
rect -194 -191 -192 -181
rect -119 -188 -117 -176
rect -109 -188 -107 -178
rect -99 -188 -97 -178
rect -33 -187 -31 -160
rect -17 -187 -15 -169
rect -7 -187 -5 -169
rect 3 -187 5 -160
rect 51 -187 53 -160
rect 67 -187 69 -169
rect 77 -187 79 -169
rect 87 -187 89 -160
rect 113 -188 115 -176
rect 123 -188 125 -178
rect 133 -188 135 -178
rect -682 -295 -680 -277
rect -675 -295 -673 -277
rect -662 -286 -660 -274
rect -353 -293 -351 -275
rect -346 -293 -344 -275
rect -333 -284 -331 -272
rect -26 -290 -24 -272
rect -19 -290 -17 -272
rect -6 -281 -4 -269
rect -776 -339 -774 -327
rect -766 -339 -764 -329
rect -756 -339 -754 -329
rect -690 -338 -688 -311
rect -674 -338 -672 -320
rect -664 -338 -662 -320
rect -654 -338 -652 -311
rect -606 -338 -604 -311
rect -590 -338 -588 -320
rect -580 -338 -578 -320
rect -570 -338 -568 -311
rect -544 -339 -542 -327
rect -534 -339 -532 -329
rect -524 -339 -522 -329
rect -447 -337 -445 -325
rect -437 -337 -435 -327
rect -427 -337 -425 -327
rect -361 -336 -359 -309
rect -345 -336 -343 -318
rect -335 -336 -333 -318
rect -325 -336 -323 -309
rect -277 -336 -275 -309
rect -261 -336 -259 -318
rect -251 -336 -249 -318
rect -241 -336 -239 -309
rect -215 -337 -213 -325
rect -205 -337 -203 -327
rect -195 -337 -193 -327
rect -120 -334 -118 -322
rect -110 -334 -108 -324
rect -100 -334 -98 -324
rect -34 -333 -32 -306
rect -18 -333 -16 -315
rect -8 -333 -6 -315
rect 2 -333 4 -306
rect 50 -333 52 -306
rect 66 -333 68 -315
rect 76 -333 78 -315
rect 86 -333 88 -306
rect 112 -334 114 -322
rect 122 -334 124 -324
rect 132 -334 134 -324
rect -683 -441 -681 -423
rect -676 -441 -674 -423
rect -663 -432 -661 -420
rect -354 -439 -352 -421
rect -347 -439 -345 -421
rect -334 -430 -332 -418
rect -27 -436 -25 -418
rect -20 -436 -18 -418
rect -7 -427 -5 -415
rect -482 -486 -480 -468
rect -472 -479 -470 -466
rect -462 -479 -460 -466
rect -389 -486 -387 -468
rect -379 -479 -377 -466
rect -369 -479 -367 -466
rect -302 -486 -300 -468
rect -292 -479 -290 -466
rect -282 -479 -280 -466
<< polycontact >>
rect -80 -50 -76 -46
rect -8 -51 -4 -47
rect 30 -51 34 -47
rect 51 -51 55 -47
rect 84 -51 88 -47
rect 105 -51 109 -47
rect 140 -51 144 -47
rect 161 -51 165 -47
rect 194 -51 198 -47
rect 215 -51 219 -47
rect -690 -114 -686 -110
rect -680 -114 -676 -110
rect -700 -122 -696 -118
rect -603 -114 -599 -110
rect -593 -114 -589 -110
rect -613 -122 -609 -118
rect -510 -114 -506 -110
rect -500 -114 -496 -110
rect -520 -122 -516 -118
rect -276 -112 -272 -108
rect -266 -112 -262 -108
rect -183 -112 -179 -108
rect -173 -112 -169 -108
rect -256 -120 -252 -116
rect -96 -112 -92 -108
rect -86 -112 -82 -108
rect -163 -120 -159 -116
rect -4 -116 0 -112
rect 34 -116 38 -112
rect 55 -116 59 -112
rect 88 -116 92 -112
rect 109 -116 113 -112
rect 144 -116 148 -112
rect 165 -116 169 -112
rect 198 -116 202 -112
rect 219 -116 223 -112
rect -76 -120 -72 -116
rect -764 -177 -760 -173
rect -703 -185 -699 -181
rect -774 -201 -770 -197
rect -619 -185 -615 -181
rect -666 -200 -662 -196
rect -656 -200 -652 -196
rect -532 -177 -528 -173
rect -435 -175 -431 -171
rect -374 -183 -370 -179
rect -755 -209 -751 -205
rect -687 -206 -683 -202
rect -582 -200 -578 -196
rect -572 -200 -568 -196
rect -542 -201 -538 -197
rect -603 -206 -599 -202
rect -445 -199 -441 -195
rect -523 -209 -519 -205
rect -290 -183 -286 -179
rect -337 -198 -333 -194
rect -327 -198 -323 -194
rect -203 -175 -199 -171
rect -108 -172 -104 -168
rect -47 -180 -43 -176
rect -426 -207 -422 -203
rect -358 -204 -354 -200
rect -253 -198 -249 -194
rect -243 -198 -239 -194
rect -213 -199 -209 -195
rect -274 -204 -270 -200
rect -118 -196 -114 -192
rect -194 -207 -190 -203
rect 37 -180 41 -176
rect -10 -195 -6 -191
rect 0 -195 4 -191
rect 124 -172 128 -168
rect -99 -204 -95 -200
rect -31 -201 -27 -197
rect 74 -195 78 -191
rect 84 -195 88 -191
rect 114 -196 118 -192
rect 53 -201 57 -197
rect 133 -204 137 -200
rect -685 -263 -681 -259
rect -673 -263 -669 -259
rect -665 -264 -661 -260
rect -356 -261 -352 -257
rect -344 -261 -340 -257
rect -675 -271 -671 -267
rect -336 -262 -332 -258
rect -29 -258 -25 -254
rect -17 -258 -13 -254
rect -346 -269 -342 -265
rect -9 -259 -5 -255
rect -19 -266 -15 -262
rect -765 -323 -761 -319
rect -704 -331 -700 -327
rect -775 -347 -771 -343
rect -620 -331 -616 -327
rect -667 -346 -663 -342
rect -657 -346 -653 -342
rect -533 -323 -529 -319
rect -436 -321 -432 -317
rect -375 -329 -371 -325
rect -756 -355 -752 -351
rect -688 -352 -684 -348
rect -583 -346 -579 -342
rect -573 -346 -569 -342
rect -543 -347 -539 -343
rect -604 -352 -600 -348
rect -446 -345 -442 -341
rect -524 -355 -520 -351
rect -291 -329 -287 -325
rect -338 -344 -334 -340
rect -328 -344 -324 -340
rect -204 -321 -200 -317
rect -109 -318 -105 -314
rect -48 -326 -44 -322
rect -427 -353 -423 -349
rect -359 -350 -355 -346
rect -254 -344 -250 -340
rect -244 -344 -240 -340
rect -214 -345 -210 -341
rect -275 -350 -271 -346
rect -119 -342 -115 -338
rect -195 -353 -191 -349
rect 36 -326 40 -322
rect -11 -341 -7 -337
rect -1 -341 3 -337
rect 123 -318 127 -314
rect -100 -350 -96 -346
rect -32 -347 -28 -343
rect 73 -341 77 -337
rect 83 -341 87 -337
rect 113 -342 117 -338
rect 52 -347 56 -343
rect 132 -350 136 -346
rect -686 -409 -682 -405
rect -674 -409 -670 -405
rect -666 -410 -662 -406
rect -357 -407 -353 -403
rect -345 -407 -341 -403
rect -676 -417 -672 -413
rect -337 -408 -333 -404
rect -30 -404 -26 -400
rect -18 -404 -14 -400
rect -347 -415 -343 -411
rect -10 -405 -6 -401
rect -20 -412 -16 -408
rect -461 -487 -457 -483
rect -481 -495 -477 -491
rect -471 -495 -467 -491
rect -368 -487 -364 -483
rect -388 -495 -384 -491
rect -378 -495 -374 -491
rect -281 -487 -277 -483
rect -301 -495 -297 -491
rect -291 -495 -287 -491
<< ndcontact >>
rect -93 -71 -89 -67
rect -59 -71 -55 -67
rect -21 -72 -17 -68
rect 13 -72 17 -68
rect 25 -71 29 -67
rect 59 -71 63 -67
rect 79 -71 83 -67
rect 113 -71 117 -67
rect 135 -71 139 -67
rect 169 -71 173 -67
rect 189 -71 193 -67
rect 223 -71 227 -67
rect -684 -88 -680 -84
rect -597 -88 -593 -84
rect -703 -98 -699 -94
rect -504 -88 -500 -84
rect -673 -100 -669 -96
rect -616 -98 -612 -94
rect -272 -86 -268 -82
rect -586 -100 -582 -96
rect -523 -98 -519 -94
rect -179 -86 -175 -82
rect -493 -100 -489 -96
rect -283 -98 -279 -94
rect -253 -96 -249 -92
rect -92 -86 -88 -82
rect -190 -98 -186 -94
rect -160 -96 -156 -92
rect -103 -98 -99 -94
rect -73 -96 -69 -92
rect -17 -95 -13 -91
rect 17 -95 21 -91
rect 29 -96 33 -92
rect 63 -96 67 -92
rect 83 -96 87 -92
rect 117 -96 121 -92
rect 139 -96 143 -92
rect 173 -96 177 -92
rect 193 -96 197 -92
rect 227 -96 231 -92
rect -781 -215 -777 -211
rect -703 -210 -699 -206
rect -619 -210 -615 -206
rect -752 -218 -748 -214
rect -689 -218 -685 -214
rect -677 -215 -673 -211
rect -667 -217 -663 -213
rect -770 -227 -766 -223
rect -605 -218 -601 -214
rect -593 -215 -589 -211
rect -583 -217 -579 -213
rect -649 -227 -645 -223
rect -549 -215 -545 -211
rect -452 -213 -448 -209
rect -374 -208 -370 -204
rect -520 -218 -516 -214
rect -290 -208 -286 -204
rect -423 -216 -419 -212
rect -360 -216 -356 -212
rect -348 -213 -344 -209
rect -338 -215 -334 -211
rect -565 -227 -561 -223
rect -538 -227 -534 -223
rect -441 -225 -437 -221
rect -276 -216 -272 -212
rect -264 -213 -260 -209
rect -254 -215 -250 -211
rect -320 -225 -316 -221
rect -220 -213 -216 -209
rect -125 -210 -121 -206
rect -47 -205 -43 -201
rect -191 -216 -187 -212
rect 37 -205 41 -201
rect -96 -213 -92 -209
rect -33 -213 -29 -209
rect -21 -210 -17 -206
rect -11 -212 -7 -208
rect -236 -225 -232 -221
rect -209 -225 -205 -221
rect -114 -222 -110 -218
rect 51 -213 55 -209
rect 63 -210 67 -206
rect 73 -212 77 -208
rect 7 -222 11 -218
rect 107 -210 111 -206
rect 136 -213 140 -209
rect 91 -222 95 -218
rect 118 -222 122 -218
rect -688 -249 -684 -245
rect -678 -249 -674 -245
rect -668 -249 -664 -245
rect -658 -249 -654 -245
rect -359 -247 -355 -243
rect -349 -247 -345 -243
rect -339 -247 -335 -243
rect -329 -247 -325 -243
rect -32 -244 -28 -240
rect -22 -244 -18 -240
rect -12 -244 -8 -240
rect -2 -244 2 -240
rect -782 -361 -778 -357
rect -704 -356 -700 -352
rect -620 -356 -616 -352
rect -753 -364 -749 -360
rect -690 -364 -686 -360
rect -678 -361 -674 -357
rect -668 -363 -664 -359
rect -771 -373 -767 -369
rect -606 -364 -602 -360
rect -594 -361 -590 -357
rect -584 -363 -580 -359
rect -650 -373 -646 -369
rect -550 -361 -546 -357
rect -453 -359 -449 -355
rect -375 -354 -371 -350
rect -521 -364 -517 -360
rect -291 -354 -287 -350
rect -424 -362 -420 -358
rect -361 -362 -357 -358
rect -349 -359 -345 -355
rect -339 -361 -335 -357
rect -566 -373 -562 -369
rect -539 -373 -535 -369
rect -442 -371 -438 -367
rect -277 -362 -273 -358
rect -265 -359 -261 -355
rect -255 -361 -251 -357
rect -321 -371 -317 -367
rect -221 -359 -217 -355
rect -126 -356 -122 -352
rect -48 -351 -44 -347
rect -192 -362 -188 -358
rect 36 -351 40 -347
rect -97 -359 -93 -355
rect -34 -359 -30 -355
rect -22 -356 -18 -352
rect -12 -358 -8 -354
rect -237 -371 -233 -367
rect -210 -371 -206 -367
rect -115 -368 -111 -364
rect 50 -359 54 -355
rect 62 -356 66 -352
rect 72 -358 76 -354
rect 6 -368 10 -364
rect 106 -356 110 -352
rect 135 -359 139 -355
rect 90 -368 94 -364
rect 117 -368 121 -364
rect -689 -395 -685 -391
rect -679 -395 -675 -391
rect -669 -395 -665 -391
rect -659 -395 -655 -391
rect -360 -393 -356 -389
rect -350 -393 -346 -389
rect -340 -393 -336 -389
rect -330 -393 -326 -389
rect -33 -390 -29 -386
rect -23 -390 -19 -386
rect -13 -390 -9 -386
rect -3 -390 1 -386
rect -488 -509 -484 -505
rect -458 -511 -454 -507
rect -395 -509 -391 -505
rect -365 -511 -361 -507
rect -308 -509 -304 -505
rect -477 -521 -473 -517
rect -278 -511 -274 -507
rect -384 -521 -380 -517
rect -297 -521 -293 -517
<< pdcontact >>
rect -104 -34 -100 -30
rect -60 -34 -54 -28
rect -21 -34 -17 -30
rect 12 -34 16 -30
rect 25 -34 29 -30
rect 42 -34 46 -30
rect 59 -34 63 -30
rect 79 -34 83 -30
rect 96 -34 100 -30
rect 113 -34 117 -30
rect 135 -34 139 -30
rect 152 -34 156 -30
rect 169 -34 173 -30
rect 189 -34 193 -30
rect 206 -34 210 -30
rect 223 -34 227 -30
rect -703 -138 -699 -134
rect -693 -131 -689 -127
rect -693 -138 -689 -134
rect -683 -136 -679 -132
rect -673 -124 -669 -120
rect -673 -131 -669 -127
rect -616 -138 -612 -134
rect -606 -131 -602 -127
rect -606 -138 -602 -134
rect -596 -136 -592 -132
rect -586 -124 -582 -120
rect -586 -131 -582 -127
rect -523 -138 -519 -134
rect -513 -131 -509 -127
rect -513 -138 -509 -134
rect -503 -136 -499 -132
rect -493 -124 -489 -120
rect -493 -131 -489 -127
rect -283 -122 -279 -118
rect -283 -129 -279 -125
rect -190 -122 -186 -118
rect -273 -134 -269 -130
rect -263 -129 -259 -125
rect -263 -136 -259 -132
rect -190 -129 -186 -125
rect -253 -136 -249 -132
rect -103 -122 -99 -118
rect -180 -134 -176 -130
rect -170 -129 -166 -125
rect -170 -136 -166 -132
rect -103 -129 -99 -125
rect -160 -136 -156 -132
rect -93 -134 -89 -130
rect -83 -129 -79 -125
rect -83 -136 -79 -132
rect -73 -136 -69 -132
rect -17 -133 -13 -129
rect 16 -133 20 -129
rect 29 -133 33 -129
rect 46 -133 50 -129
rect 63 -133 67 -129
rect 83 -133 87 -129
rect 100 -133 104 -129
rect 117 -133 121 -129
rect 139 -133 143 -129
rect 156 -133 160 -129
rect 173 -133 177 -129
rect 193 -133 197 -129
rect 210 -133 214 -129
rect 227 -133 231 -129
rect -781 -192 -777 -188
rect -771 -192 -767 -188
rect -761 -192 -757 -188
rect -751 -188 -747 -184
rect -695 -191 -691 -187
rect -685 -170 -681 -166
rect -685 -177 -681 -173
rect -669 -191 -665 -187
rect -659 -184 -655 -180
rect -649 -176 -645 -172
rect -611 -191 -607 -187
rect -601 -170 -597 -166
rect -601 -177 -597 -173
rect -585 -191 -581 -187
rect -575 -184 -571 -180
rect -565 -176 -561 -172
rect -549 -192 -545 -188
rect -539 -192 -535 -188
rect -529 -192 -525 -188
rect -519 -188 -515 -184
rect -452 -190 -448 -186
rect -442 -190 -438 -186
rect -432 -190 -428 -186
rect -422 -186 -418 -182
rect -366 -189 -362 -185
rect -356 -168 -352 -164
rect -356 -175 -352 -171
rect -340 -189 -336 -185
rect -330 -182 -326 -178
rect -320 -174 -316 -170
rect -282 -189 -278 -185
rect -272 -168 -268 -164
rect -272 -175 -268 -171
rect -256 -189 -252 -185
rect -246 -182 -242 -178
rect -236 -174 -232 -170
rect -220 -190 -216 -186
rect -210 -190 -206 -186
rect -200 -190 -196 -186
rect -190 -186 -186 -182
rect -125 -187 -121 -183
rect -115 -187 -111 -183
rect -105 -187 -101 -183
rect -95 -183 -91 -179
rect -39 -186 -35 -182
rect -29 -165 -25 -161
rect -29 -172 -25 -168
rect -13 -186 -9 -182
rect -3 -179 1 -175
rect 7 -171 11 -167
rect 45 -186 49 -182
rect 55 -165 59 -161
rect 55 -172 59 -168
rect 71 -186 75 -182
rect 81 -179 85 -175
rect 91 -171 95 -167
rect 107 -187 111 -183
rect 117 -187 121 -183
rect 127 -187 131 -183
rect 137 -183 141 -179
rect -688 -287 -684 -283
rect -658 -285 -654 -281
rect -359 -285 -355 -281
rect -670 -294 -666 -290
rect -329 -283 -325 -279
rect -32 -282 -28 -278
rect -341 -292 -337 -288
rect -2 -280 2 -276
rect -14 -289 -10 -285
rect -782 -338 -778 -334
rect -772 -338 -768 -334
rect -762 -338 -758 -334
rect -752 -334 -748 -330
rect -696 -337 -692 -333
rect -686 -316 -682 -312
rect -686 -323 -682 -319
rect -670 -337 -666 -333
rect -660 -330 -656 -326
rect -650 -322 -646 -318
rect -612 -337 -608 -333
rect -602 -316 -598 -312
rect -602 -323 -598 -319
rect -586 -337 -582 -333
rect -576 -330 -572 -326
rect -566 -322 -562 -318
rect -550 -338 -546 -334
rect -540 -338 -536 -334
rect -530 -338 -526 -334
rect -520 -334 -516 -330
rect -453 -336 -449 -332
rect -443 -336 -439 -332
rect -433 -336 -429 -332
rect -423 -332 -419 -328
rect -367 -335 -363 -331
rect -357 -314 -353 -310
rect -357 -321 -353 -317
rect -341 -335 -337 -331
rect -331 -328 -327 -324
rect -321 -320 -317 -316
rect -283 -335 -279 -331
rect -273 -314 -269 -310
rect -273 -321 -269 -317
rect -257 -335 -253 -331
rect -247 -328 -243 -324
rect -237 -320 -233 -316
rect -221 -336 -217 -332
rect -211 -336 -207 -332
rect -201 -336 -197 -332
rect -191 -332 -187 -328
rect -126 -333 -122 -329
rect -116 -333 -112 -329
rect -106 -333 -102 -329
rect -96 -329 -92 -325
rect -40 -332 -36 -328
rect -30 -311 -26 -307
rect -30 -318 -26 -314
rect -14 -332 -10 -328
rect -4 -325 0 -321
rect 6 -317 10 -313
rect 44 -332 48 -328
rect 54 -311 58 -307
rect 54 -318 58 -314
rect 70 -332 74 -328
rect 80 -325 84 -321
rect 90 -317 94 -313
rect 106 -333 110 -329
rect 116 -333 120 -329
rect 126 -333 130 -329
rect 136 -329 140 -325
rect -689 -433 -685 -429
rect -659 -431 -655 -427
rect -360 -431 -356 -427
rect -671 -440 -667 -436
rect -330 -429 -326 -425
rect -33 -428 -29 -424
rect -342 -438 -338 -434
rect -3 -426 1 -422
rect -15 -435 -11 -431
rect -488 -478 -484 -474
rect -488 -485 -484 -481
rect -478 -473 -474 -469
rect -468 -471 -464 -467
rect -468 -478 -464 -474
rect -458 -471 -454 -467
rect -395 -478 -391 -474
rect -395 -485 -391 -481
rect -385 -473 -381 -469
rect -375 -471 -371 -467
rect -375 -478 -371 -474
rect -365 -471 -361 -467
rect -308 -478 -304 -474
rect -308 -485 -304 -481
rect -298 -473 -294 -469
rect -288 -471 -284 -467
rect -288 -478 -284 -474
rect -278 -471 -274 -467
<< m2contact >>
rect -73 -49 -69 -45
rect -1 -50 3 -46
rect -58 -59 -54 -55
rect 24 -50 28 -46
rect 46 -50 50 -46
rect 66 -42 70 -38
rect 76 -50 80 -46
rect -344 -72 -339 -66
rect 14 -60 18 -56
rect 100 -59 104 -55
rect 133 -50 137 -46
rect 169 -47 173 -43
rect 132 -58 136 -54
rect 149 -55 153 -51
rect 159 -57 163 -53
rect 122 -65 126 -61
rect 208 -49 212 -45
rect 222 -56 226 -52
rect 191 -64 195 -60
rect -708 -81 -703 -76
rect -786 -99 -781 -93
rect -708 -105 -704 -101
rect -716 -131 -711 -126
rect -620 -105 -616 -101
rect -624 -131 -620 -127
rect -527 -105 -523 -101
rect -479 -100 -475 -96
rect -303 -100 -298 -95
rect -575 -132 -571 -128
rect -531 -131 -527 -127
rect -345 -111 -340 -106
rect -249 -103 -245 -99
rect -479 -123 -475 -119
rect -302 -123 -297 -118
rect -245 -129 -241 -125
rect -479 -140 -475 -136
rect -301 -140 -297 -136
rect -214 -130 -210 -125
rect -156 -104 -152 -100
rect -69 -104 -65 -100
rect -45 -102 -41 -98
rect 10 -100 14 -96
rect 18 -107 22 -103
rect -152 -129 -148 -125
rect -139 -127 -135 -123
rect -586 -157 -582 -153
rect -549 -156 -544 -152
rect -238 -151 -233 -146
rect -203 -151 -199 -146
rect -140 -151 -136 -147
rect -126 -152 -122 -148
rect -116 -127 -112 -123
rect 3 -117 7 -113
rect -64 -129 -59 -125
rect 74 -100 78 -96
rect 28 -117 32 -113
rect 50 -117 54 -113
rect 80 -117 84 -113
rect 104 -108 108 -104
rect 96 -117 100 -113
rect 136 -109 140 -105
rect 72 -125 76 -121
rect 163 -110 167 -106
rect 137 -117 141 -113
rect 195 -103 199 -99
rect 226 -111 230 -107
rect 173 -120 177 -116
rect 212 -118 216 -114
rect -116 -151 -112 -147
rect -758 -177 -754 -173
rect -615 -177 -611 -173
rect -782 -205 -778 -201
rect -750 -203 -746 -199
rect -713 -203 -709 -199
rect -693 -204 -689 -200
rect -646 -204 -642 -200
rect -609 -204 -605 -200
rect -526 -177 -522 -173
rect -557 -220 -553 -216
rect -518 -202 -514 -198
rect -801 -231 -797 -227
rect -516 -230 -510 -224
rect -689 -272 -685 -268
rect -698 -280 -694 -276
rect -496 -254 -492 -250
rect -429 -175 -425 -171
rect -286 -175 -282 -171
rect -453 -203 -449 -199
rect -421 -201 -417 -197
rect -384 -201 -380 -197
rect -364 -202 -360 -198
rect -229 -182 -225 -178
rect -317 -202 -313 -198
rect -280 -202 -276 -198
rect -197 -175 -193 -171
rect -228 -218 -224 -214
rect -189 -200 -185 -196
rect -476 -231 -469 -224
rect -189 -228 -183 -222
rect -471 -254 -467 -250
rect -399 -254 -395 -250
rect -360 -270 -356 -266
rect -369 -278 -365 -274
rect -177 -257 -173 -253
rect -102 -172 -98 -168
rect 41 -172 45 -168
rect -67 -182 -63 -178
rect -126 -200 -122 -196
rect -94 -198 -90 -194
rect -57 -198 -53 -194
rect -37 -199 -33 -195
rect 18 -180 22 -176
rect 10 -199 14 -195
rect -66 -215 -62 -211
rect 19 -215 23 -211
rect 96 -179 101 -175
rect 47 -199 51 -195
rect 130 -172 134 -168
rect 99 -215 103 -211
rect 138 -197 142 -193
rect -149 -229 -142 -222
rect -65 -245 -60 -240
rect -145 -257 -141 -253
rect -74 -257 -70 -253
rect -516 -302 -511 -298
rect -496 -303 -491 -298
rect -52 -252 -48 -248
rect -33 -267 -29 -263
rect -42 -275 -38 -271
rect 11 -252 15 -248
rect 19 -258 23 -253
rect -52 -283 -48 -279
rect -64 -289 -60 -285
rect 18 -293 23 -286
rect -759 -323 -755 -319
rect -783 -351 -779 -347
rect -751 -349 -747 -345
rect -714 -349 -710 -345
rect -694 -350 -690 -346
rect -647 -350 -643 -346
rect -616 -323 -612 -319
rect -610 -350 -606 -346
rect -633 -366 -629 -362
rect -527 -323 -523 -319
rect -558 -366 -554 -362
rect -519 -348 -515 -344
rect -516 -376 -508 -369
rect -567 -386 -563 -382
rect -690 -418 -686 -414
rect -699 -426 -695 -422
rect -572 -405 -566 -399
rect -543 -405 -538 -400
rect -518 -405 -513 -400
rect -497 -405 -492 -400
rect -430 -321 -426 -317
rect -287 -321 -283 -317
rect -394 -340 -390 -336
rect -454 -349 -450 -345
rect -422 -347 -418 -343
rect -385 -347 -381 -343
rect -365 -348 -361 -344
rect -318 -348 -314 -344
rect -394 -364 -390 -360
rect -281 -348 -277 -344
rect -198 -321 -194 -317
rect -229 -364 -225 -360
rect -190 -346 -186 -342
rect -479 -376 -474 -371
rect -189 -375 -185 -371
rect -394 -390 -390 -386
rect -394 -408 -390 -404
rect -361 -416 -357 -412
rect -370 -424 -366 -420
rect -304 -398 -298 -393
rect -216 -398 -211 -393
rect -103 -318 -99 -314
rect 40 -318 44 -314
rect -127 -346 -123 -342
rect -95 -344 -91 -340
rect -58 -344 -54 -340
rect -38 -345 -34 -341
rect 9 -345 13 -341
rect 46 -345 50 -341
rect 129 -318 133 -314
rect 98 -361 102 -357
rect 137 -343 141 -339
rect -149 -375 -145 -371
rect -91 -384 -87 -380
rect -152 -398 -147 -393
rect -118 -398 -113 -393
rect -321 -431 -316 -426
rect -422 -438 -418 -434
rect -34 -413 -30 -409
rect -43 -421 -39 -417
rect 14 -396 20 -391
rect -91 -425 -87 -421
rect -422 -467 -418 -463
rect -450 -504 -445 -499
rect -430 -515 -426 -511
rect -320 -475 -316 -470
rect -353 -487 -349 -482
rect -357 -504 -352 -499
rect -264 -487 -260 -483
rect -272 -504 -267 -499
rect -506 -526 -499 -519
<< m3contact >>
rect -320 -155 -316 -151
rect -301 -176 -297 -172
<< psubstratepcontact >>
rect -674 -88 -670 -84
rect -587 -88 -583 -84
rect -494 -88 -490 -84
rect -282 -86 -278 -82
rect -189 -86 -185 -82
rect -102 -86 -98 -82
rect -780 -227 -776 -223
rect -702 -227 -698 -223
rect -618 -227 -614 -223
rect -548 -227 -544 -223
rect -451 -225 -447 -221
rect -373 -225 -369 -221
rect -289 -225 -285 -221
rect -219 -225 -215 -221
rect -124 -222 -120 -218
rect -46 -222 -42 -218
rect 38 -222 42 -218
rect 108 -222 112 -218
rect -687 -237 -683 -233
rect -659 -237 -655 -233
rect -358 -235 -354 -231
rect -330 -235 -326 -231
rect -31 -232 -27 -228
rect -3 -232 1 -228
rect -781 -373 -777 -369
rect -703 -373 -699 -369
rect -619 -373 -615 -369
rect -549 -373 -545 -369
rect -452 -371 -448 -367
rect -374 -371 -370 -367
rect -290 -371 -286 -367
rect -220 -371 -216 -367
rect -125 -368 -121 -364
rect -47 -368 -43 -364
rect 37 -368 41 -364
rect 107 -368 111 -364
rect -688 -383 -684 -379
rect -660 -383 -656 -379
rect -359 -381 -355 -377
rect -331 -381 -327 -377
rect -32 -378 -28 -374
rect -4 -378 0 -374
rect -487 -521 -483 -517
rect -394 -521 -390 -517
rect -307 -521 -303 -517
<< nsubstratencontact >>
rect 52 -20 56 -16
rect 106 -20 110 -16
rect 162 -20 166 -16
rect 216 -20 220 -16
rect -674 -148 -670 -144
rect -587 -148 -583 -144
rect -494 -148 -490 -144
rect -282 -146 -278 -142
rect -189 -146 -185 -142
rect -102 -146 -98 -142
rect 56 -147 60 -143
rect 110 -147 114 -143
rect 166 -147 170 -143
rect 220 -147 224 -143
rect -780 -167 -776 -163
rect -766 -167 -762 -163
rect -752 -167 -748 -163
rect -669 -167 -665 -163
rect -585 -167 -581 -163
rect -548 -167 -544 -163
rect -534 -167 -530 -163
rect -520 -167 -516 -163
rect -451 -165 -447 -161
rect -437 -165 -433 -161
rect -423 -165 -419 -161
rect -340 -165 -336 -161
rect -256 -165 -252 -161
rect -219 -165 -215 -161
rect -205 -165 -201 -161
rect -191 -165 -187 -161
rect -124 -162 -120 -158
rect -110 -162 -106 -158
rect -96 -162 -92 -158
rect -13 -162 -9 -158
rect 71 -162 75 -158
rect 108 -162 112 -158
rect 122 -162 126 -158
rect 136 -162 140 -158
rect -659 -297 -655 -293
rect -330 -295 -326 -291
rect -3 -292 1 -288
rect -781 -313 -777 -309
rect -767 -313 -763 -309
rect -753 -313 -749 -309
rect -670 -313 -666 -309
rect -586 -313 -582 -309
rect -549 -313 -545 -309
rect -535 -313 -531 -309
rect -521 -313 -517 -309
rect -452 -311 -448 -307
rect -438 -311 -434 -307
rect -424 -311 -420 -307
rect -341 -311 -337 -307
rect -257 -311 -253 -307
rect -220 -311 -216 -307
rect -206 -311 -202 -307
rect -192 -311 -188 -307
rect -125 -308 -121 -304
rect -111 -308 -107 -304
rect -97 -308 -93 -304
rect -14 -308 -10 -304
rect 70 -308 74 -304
rect 107 -308 111 -304
rect 121 -308 125 -304
rect 135 -308 139 -304
rect -660 -443 -656 -439
rect -331 -441 -327 -437
rect -4 -438 0 -434
rect -487 -461 -483 -457
rect -394 -461 -390 -457
rect -307 -461 -303 -457
<< psubstratepdiff >>
rect -283 -82 -277 -81
rect -675 -84 -669 -83
rect -675 -88 -674 -84
rect -670 -88 -669 -84
rect -675 -89 -669 -88
rect -588 -84 -582 -83
rect -588 -88 -587 -84
rect -583 -88 -582 -84
rect -588 -89 -582 -88
rect -495 -84 -489 -83
rect -495 -88 -494 -84
rect -490 -88 -489 -84
rect -283 -86 -282 -82
rect -278 -86 -277 -82
rect -283 -87 -277 -86
rect -190 -82 -184 -81
rect -190 -86 -189 -82
rect -185 -86 -184 -82
rect -495 -89 -489 -88
rect -190 -87 -184 -86
rect -103 -82 -97 -81
rect -103 -86 -102 -82
rect -98 -86 -97 -82
rect -103 -87 -97 -86
rect -781 -223 -775 -222
rect -781 -227 -780 -223
rect -776 -227 -775 -223
rect -781 -228 -775 -227
rect -703 -223 -697 -222
rect -703 -227 -702 -223
rect -698 -227 -697 -223
rect -703 -228 -697 -227
rect -619 -223 -613 -222
rect -619 -227 -618 -223
rect -614 -227 -613 -223
rect -619 -228 -613 -227
rect -452 -221 -446 -220
rect -549 -223 -543 -222
rect -549 -227 -548 -223
rect -544 -227 -543 -223
rect -549 -228 -543 -227
rect -452 -225 -451 -221
rect -447 -225 -446 -221
rect -452 -226 -446 -225
rect -374 -221 -368 -220
rect -374 -225 -373 -221
rect -369 -225 -368 -221
rect -374 -226 -368 -225
rect -290 -221 -284 -220
rect -290 -225 -289 -221
rect -285 -225 -284 -221
rect -290 -226 -284 -225
rect -125 -218 -119 -217
rect -220 -221 -214 -220
rect -220 -225 -219 -221
rect -215 -225 -214 -221
rect -220 -226 -214 -225
rect -125 -222 -124 -218
rect -120 -222 -119 -218
rect -125 -223 -119 -222
rect -47 -218 -41 -217
rect -47 -222 -46 -218
rect -42 -222 -41 -218
rect -47 -223 -41 -222
rect 37 -218 43 -217
rect 37 -222 38 -218
rect 42 -222 43 -218
rect 37 -223 43 -222
rect 107 -218 113 -217
rect 107 -222 108 -218
rect 112 -222 113 -218
rect 107 -223 113 -222
rect -32 -228 2 -227
rect -359 -231 -325 -230
rect -688 -233 -654 -232
rect -688 -237 -687 -233
rect -683 -237 -659 -233
rect -655 -237 -654 -233
rect -359 -235 -358 -231
rect -354 -235 -330 -231
rect -326 -235 -325 -231
rect -32 -232 -31 -228
rect -27 -232 -3 -228
rect 1 -232 2 -228
rect -32 -233 2 -232
rect -359 -236 -325 -235
rect -688 -238 -654 -237
rect -782 -369 -776 -368
rect -782 -373 -781 -369
rect -777 -373 -776 -369
rect -782 -374 -776 -373
rect -704 -369 -698 -368
rect -704 -373 -703 -369
rect -699 -373 -698 -369
rect -704 -374 -698 -373
rect -620 -369 -614 -368
rect -620 -373 -619 -369
rect -615 -373 -614 -369
rect -620 -374 -614 -373
rect -453 -367 -447 -366
rect -550 -369 -544 -368
rect -550 -373 -549 -369
rect -545 -373 -544 -369
rect -550 -374 -544 -373
rect -453 -371 -452 -367
rect -448 -371 -447 -367
rect -453 -372 -447 -371
rect -375 -367 -369 -366
rect -375 -371 -374 -367
rect -370 -371 -369 -367
rect -375 -372 -369 -371
rect -291 -367 -285 -366
rect -291 -371 -290 -367
rect -286 -371 -285 -367
rect -291 -372 -285 -371
rect -126 -364 -120 -363
rect -221 -367 -215 -366
rect -221 -371 -220 -367
rect -216 -371 -215 -367
rect -221 -372 -215 -371
rect -126 -368 -125 -364
rect -121 -368 -120 -364
rect -126 -369 -120 -368
rect -48 -364 -42 -363
rect -48 -368 -47 -364
rect -43 -368 -42 -364
rect -48 -369 -42 -368
rect 36 -364 42 -363
rect 36 -368 37 -364
rect 41 -368 42 -364
rect 36 -369 42 -368
rect 106 -364 112 -363
rect 106 -368 107 -364
rect 111 -368 112 -364
rect 106 -369 112 -368
rect -33 -374 1 -373
rect -360 -377 -326 -376
rect -689 -379 -655 -378
rect -689 -383 -688 -379
rect -684 -383 -660 -379
rect -656 -383 -655 -379
rect -360 -381 -359 -377
rect -355 -381 -331 -377
rect -327 -381 -326 -377
rect -33 -378 -32 -374
rect -28 -378 -4 -374
rect 0 -378 1 -374
rect -33 -379 1 -378
rect -360 -382 -326 -381
rect -689 -384 -655 -383
rect -488 -517 -482 -516
rect -488 -521 -487 -517
rect -483 -521 -482 -517
rect -488 -522 -482 -521
rect -395 -517 -389 -516
rect -395 -521 -394 -517
rect -390 -521 -389 -517
rect -395 -522 -389 -521
rect -308 -517 -302 -516
rect -308 -521 -307 -517
rect -303 -521 -302 -517
rect -308 -522 -302 -521
<< nsubstratendiff >>
rect -675 -144 -669 -143
rect -588 -144 -582 -143
rect -283 -142 -277 -141
rect -190 -142 -184 -141
rect -103 -142 -97 -141
rect -495 -144 -489 -143
rect -675 -148 -674 -144
rect -670 -148 -669 -144
rect -675 -149 -669 -148
rect -588 -148 -587 -144
rect -583 -148 -582 -144
rect -588 -149 -582 -148
rect -495 -148 -494 -144
rect -490 -148 -489 -144
rect -283 -146 -282 -142
rect -278 -146 -277 -142
rect -283 -147 -277 -146
rect -190 -146 -189 -142
rect -185 -146 -184 -142
rect -190 -147 -184 -146
rect -103 -146 -102 -142
rect -98 -146 -97 -142
rect -103 -147 -97 -146
rect -495 -149 -489 -148
rect -452 -161 -418 -160
rect -781 -163 -747 -162
rect -781 -167 -780 -163
rect -776 -167 -766 -163
rect -762 -167 -752 -163
rect -748 -167 -747 -163
rect -670 -163 -664 -162
rect -781 -168 -747 -167
rect -670 -167 -669 -163
rect -665 -167 -664 -163
rect -586 -163 -580 -162
rect -670 -168 -664 -167
rect -586 -167 -585 -163
rect -581 -167 -580 -163
rect -549 -163 -515 -162
rect -586 -168 -580 -167
rect -549 -167 -548 -163
rect -544 -167 -534 -163
rect -530 -167 -520 -163
rect -516 -167 -515 -163
rect -452 -165 -451 -161
rect -447 -165 -437 -161
rect -433 -165 -423 -161
rect -419 -165 -418 -161
rect -341 -161 -335 -160
rect -452 -166 -418 -165
rect -549 -168 -515 -167
rect -341 -165 -340 -161
rect -336 -165 -335 -161
rect -257 -161 -251 -160
rect -341 -166 -335 -165
rect -257 -165 -256 -161
rect -252 -165 -251 -161
rect -220 -161 -186 -160
rect -257 -166 -251 -165
rect -220 -165 -219 -161
rect -215 -165 -205 -161
rect -201 -165 -191 -161
rect -187 -165 -186 -161
rect -125 -162 -124 -158
rect -120 -162 -110 -158
rect -106 -162 -96 -158
rect -92 -162 -91 -158
rect -14 -158 -8 -157
rect -125 -163 -91 -162
rect -220 -166 -186 -165
rect -14 -162 -13 -158
rect -9 -162 -8 -158
rect 70 -158 76 -157
rect -14 -163 -8 -162
rect 70 -162 71 -158
rect 75 -162 76 -158
rect 107 -158 141 -157
rect 70 -163 76 -162
rect 107 -162 108 -158
rect 112 -162 122 -158
rect 126 -162 136 -158
rect 140 -162 141 -158
rect 107 -163 141 -162
rect -660 -293 -654 -292
rect -4 -288 2 -287
rect -331 -291 -325 -290
rect -660 -297 -659 -293
rect -655 -297 -654 -293
rect -331 -295 -330 -291
rect -326 -295 -325 -291
rect -4 -292 -3 -288
rect 1 -292 2 -288
rect -4 -293 2 -292
rect -331 -296 -325 -295
rect -660 -298 -654 -297
rect -126 -304 -92 -303
rect -453 -307 -419 -306
rect -782 -309 -748 -308
rect -782 -313 -781 -309
rect -777 -313 -767 -309
rect -763 -313 -753 -309
rect -749 -313 -748 -309
rect -671 -309 -665 -308
rect -782 -314 -748 -313
rect -671 -313 -670 -309
rect -666 -313 -665 -309
rect -587 -309 -581 -308
rect -671 -314 -665 -313
rect -587 -313 -586 -309
rect -582 -313 -581 -309
rect -550 -309 -516 -308
rect -587 -314 -581 -313
rect -550 -313 -549 -309
rect -545 -313 -535 -309
rect -531 -313 -521 -309
rect -517 -313 -516 -309
rect -453 -311 -452 -307
rect -448 -311 -438 -307
rect -434 -311 -424 -307
rect -420 -311 -419 -307
rect -342 -307 -336 -306
rect -453 -312 -419 -311
rect -550 -314 -516 -313
rect -342 -311 -341 -307
rect -337 -311 -336 -307
rect -258 -307 -252 -306
rect -342 -312 -336 -311
rect -258 -311 -257 -307
rect -253 -311 -252 -307
rect -221 -307 -187 -306
rect -258 -312 -252 -311
rect -221 -311 -220 -307
rect -216 -311 -206 -307
rect -202 -311 -192 -307
rect -188 -311 -187 -307
rect -126 -308 -125 -304
rect -121 -308 -111 -304
rect -107 -308 -97 -304
rect -93 -308 -92 -304
rect -15 -304 -9 -303
rect -126 -309 -92 -308
rect -221 -312 -187 -311
rect -15 -308 -14 -304
rect -10 -308 -9 -304
rect 69 -304 75 -303
rect -15 -309 -9 -308
rect 69 -308 70 -304
rect 74 -308 75 -304
rect 106 -304 140 -303
rect 69 -309 75 -308
rect 106 -308 107 -304
rect 111 -308 121 -304
rect 125 -308 135 -304
rect 139 -308 140 -304
rect 106 -309 140 -308
rect -661 -439 -655 -438
rect -5 -434 1 -433
rect -332 -437 -326 -436
rect -661 -443 -660 -439
rect -656 -443 -655 -439
rect -332 -441 -331 -437
rect -327 -441 -326 -437
rect -5 -438 -4 -434
rect 0 -438 1 -434
rect -5 -439 1 -438
rect -332 -442 -326 -441
rect -661 -444 -655 -443
rect -488 -457 -482 -456
rect -488 -461 -487 -457
rect -483 -461 -482 -457
rect -395 -457 -389 -456
rect -395 -461 -394 -457
rect -390 -461 -389 -457
rect -308 -457 -302 -456
rect -308 -461 -307 -457
rect -303 -461 -302 -457
rect -488 -462 -482 -461
rect -395 -462 -389 -461
rect -308 -462 -302 -461
<< pad >>
rect -647 -154 -643 -150
<< labels >>
rlabel metal1 -342 -231 -342 -231 2 vss
rlabel metal1 -108 -222 -108 -222 6 vss
rlabel metal1 124 -158 124 -158 6 vdd
rlabel metal1 -15 -228 -15 -228 2 vss
rlabel metal1 -15 -292 -15 -292 2 vdd
rlabel metal1 -16 -438 -16 -438 2 vdd
rlabel metal1 -16 -374 -16 -374 2 vss
rlabel metal1 123 -368 123 -368 6 vss
rlabel metal1 123 -304 123 -304 6 vdd
rlabel metal1 -109 -304 -109 -304 6 vdd
rlabel metal1 -109 -368 -109 -368 6 vss
rlabel metal1 -19 -304 -19 -304 6 vdd
rlabel metal1 -343 -377 -343 -377 2 vss
rlabel metal1 -204 -371 -204 -371 6 vss
rlabel metal1 -204 -307 -204 -307 6 vdd
rlabel metal1 -436 -307 -436 -307 6 vdd
rlabel metal1 -436 -371 -436 -371 6 vss
rlabel metal1 -262 -307 -262 -307 6 vdd
rlabel metal1 -262 -371 -262 -371 6 vss
rlabel metal1 -672 -443 -672 -443 2 vdd
rlabel metal1 -765 -309 -765 -309 6 vdd
rlabel metal1 -765 -373 -765 -373 6 vss
rlabel metal1 -591 -309 -591 -309 6 vdd
rlabel metal1 -591 -373 -591 -373 6 vss
rlabel m2contact -706 -104 -706 -104 1 q0_M1
rlabel metal1 -670 -112 -670 -112 1 q0b2_M1
rlabel metal1 -498 -105 -498 -105 1 q0b0_n_M1
rlabel metal1 -378 -99 -378 -99 1 b2_M1
rlabel metal1 -377 -120 -377 -120 1 b1_M1
rlabel metal1 -377 -139 -377 -139 1 b0_M1
rlabel metal1 -283 -101 -283 -101 1 q1b0_M1
rlabel metal1 -181 -94 -181 -94 1 q1b1_M1
rlabel metal1 -181 -116 -181 -116 1 q1b1_n_M1
rlabel metal1 -103 -105 -103 -105 1 q1b2_M1
rlabel metal1 -94 -105 -94 -105 1 q1b2_n_M1
rlabel m2contact -67 -102 -67 -102 1 q1_M1
rlabel metal1 122 -194 122 -194 1 zc1_n_3_M1
rlabel metal1 108 -194 108 -194 1 c1_3_M1
rlabel metal1 94 -190 94 -190 1 s_fa3_M1
rlabel metal1 71 -172 71 -172 1 cn_3_M1
rlabel ntransistor 87 -207 87 -207 1 s_fa3_n_M1
rlabel metal1 10 -190 10 -190 1 so_3_M1
rlabel metal1 -2 -169 -2 -169 1 bn3_M1
rlabel ptransistor -6 -185 -6 -185 1 an3_M1
rlabel metal1 -103 -190 -103 -190 1 co_n3_M1
rlabel metal1 -116 -210 -116 -210 1 co_3_M1
rlabel metal1 -219 -197 -219 -197 1 c1_2_M1
rlabel metal1 -205 -197 -205 -197 1 zc1_2_n_M1
rlabel ntransistor -240 -210 -240 -210 1 son_2_M1
rlabel pdcontact -243 -180 -243 -180 1 s_fa2_M1
rlabel metal1 -255 -197 -255 -197 1 cn2_M1
rlabel metal1 -317 -193 -317 -193 1 so_2_M1
rlabel polycontact -327 -197 -327 -197 1 an_2_M1
rlabel polycontact -333 -196 -333 -196 1 bn_2_M1
rlabel metal1 -430 -194 -430 -194 1 co_n2_M1
rlabel metal1 -443 -213 -443 -213 1 co_2_M1
rlabel metal1 -534 -199 -534 -199 1 zc1_n1_M1
rlabel metal1 -548 -199 -548 -199 1 c1_1_M1
rlabel metal1 -562 -195 -562 -195 1 a1_M1
rlabel ntransistor -569 -212 -569 -212 1 a1_n_M1
rlabel ntransistor -653 -211 -653 -211 1 an_1_M1
rlabel metal1 -646 -195 -646 -195 1 so_1_M1
rlabel metal1 -658 -174 -658 -174 1 bn_1_M1
rlabel metal1 -759 -195 -759 -195 1 co_n1_M1
rlabel metal1 -772 -215 -772 -215 1 co_1_M1
rlabel metal1 -663 -267 -663 -267 1 c_fa1_n_M1
rlabel metal1 -655 -267 -655 -267 1 c_fa1_M1
rlabel metal1 -334 -263 -334 -263 1 c_fa_n_M1
rlabel metal1 -326 -259 -326 -259 1 c_fa2_M1
rlabel metal1 -7 -260 -7 -260 1 c_fa3_n_M1
rlabel metal1 1 -256 1 -256 1 c_fa3_M1
rlabel metal1 121 -340 121 -340 1 zc1_6_n_M1
rlabel metal1 107 -340 107 -340 1 c1_6_M1
rlabel ntransistor 86 -353 86 -353 1 s_fa_6_n_M1
rlabel metal1 93 -336 93 -336 1 a2_M1
rlabel metal1 69 -319 69 -319 1 cn_6_M1
rlabel metal1 9 -336 9 -336 1 so_6_M1
rlabel ptransistor -7 -331 -7 -331 1 an_6_M1
rlabel metal1 -46 -342 -46 -342 1 bn_6_M1
rlabel metal1 -104 -336 -104 -336 1 co_n_6_M1
rlabel metal1 -117 -356 -117 -356 1 co_6_M1
rlabel metal1 -206 -343 -206 -343 1 zc1_n_5_M1
rlabel metal1 -220 -343 -220 -343 1 c1_5_M1
rlabel metal1 -258 -323 -258 -323 1 cn_5_M1
rlabel metal1 -234 -339 -234 -339 1 a3_M1
rlabel ntransistor -241 -356 -241 -356 1 s_fa5_n_M1
rlabel metal1 -330 -318 -330 -318 1 bn_5_M1
rlabel ptransistor -334 -334 -334 -334 1 an_5_M1
rlabel metal1 -318 -339 -318 -339 1 so_5_M1
rlabel metal1 -431 -339 -431 -339 1 co_5__M1
rlabel metal1 -535 -345 -535 -345 1 zc1_4_M1
rlabel metal1 -549 -345 -549 -345 1 c1_4_M1
rlabel metal1 -563 -341 -563 -341 1 a4_M1
rlabel ntransistor -570 -358 -570 -358 1 s_fa4_n_M1
rlabel metal1 -587 -325 -587 -325 1 cn_1_M1
rlabel metal1 -670 -326 -670 -326 1 bn4_M1
rlabel ptransistor -663 -336 -663 -336 1 an4_M1
rlabel metal1 -647 -341 -647 -341 1 so_4_M1
rlabel metal1 -760 -341 -760 -341 1 co_n4_M1
rlabel metal1 -773 -361 -773 -361 1 co_4_M1
rlabel metal1 -664 -411 -664 -411 1 a5_n_M1
rlabel metal1 -656 -407 -656 -407 1 a5_M1
rlabel metal1 -327 -405 -327 -405 1 c_fa5_M1
rlabel metal1 -335 -409 -335 -409 1 c_fa5_n_M1
rlabel metal1 -8 -406 -8 -406 1 c_fa6_n_M1
rlabel metal1 0 -402 0 -402 1 c_fa6_M1
rlabel metal1 -307 -499 -307 -499 1 q2b0_M1
rlabel metal1 -298 -500 -298 -500 1 q2b0_n_M1
rlabel m2contact -270 -501 -270 -501 1 q2_M1
rlabel metal1 -395 -499 -395 -499 1 q2b1_M1
rlabel metal1 -386 -499 -386 -499 1 q2b1_n_M1
rlabel metal1 -465 -510 -465 -510 1 q2b2_n_M1
rlabel metal1 -487 -511 -487 -511 1 q2b2_M1
rlabel metal1 -678 -108 -678 -108 1 q0b2_n_M1
rlabel metal1 -583 -108 -583 -108 1 q0b1_M1
rlabel metal1 -274 -115 -274 -115 1 q1b0_n_M1
rlabel metal1 -591 -107 -591 -107 1 q0b1_n_M1
rlabel metal1 -491 -106 -491 -106 1 a0_M1
rlabel metal1 18 -110 18 -110 1 n6
rlabel ndiffusion 46 -94 46 -94 1 n7
rlabel metal1 65 -111 65 -111 1 out_n7
rlabel metal1 120 -107 120 -107 1 out_n8
rlabel ndiffusion 102 -94 102 -94 1 n8
rlabel ndiffusion 158 -94 158 -94 1 n9
rlabel ndiffusion 212 -94 212 -94 1 n10
rlabel m2contact 225 -53 225 -53 1 q_l1_bar
rlabel polycontact 36 -114 36 -114 1 q_l1
rlabel m2contact -57 -57 -57 -57 1 en_bar
rlabel metal1 212 -84 212 -84 5 gnd
rlabel metal1 212 -153 212 -153 1 vdd
rlabel m2contact 229 -110 229 -110 7 q_bar
rlabel m2contact 175 -118 175 -118 5 q
rlabel metal1 61 -52 61 -52 1 out_n1
rlabel metal1 116 -56 116 -56 1 out_n2
rlabel ndiffusion 208 -69 208 -69 1 n4
rlabel ndiffusion 154 -69 154 -69 1 n3
rlabel ndiffusion 98 -69 98 -69 1 n2
rlabel ndiffusion 42 -69 42 -69 1 n1
rlabel polycontact 53 -49 53 -49 1 en
rlabel metal1 14 -50 14 -50 1 D_bar
rlabel polycontact 32 -49 32 -49 1 D
rlabel metal1 208 -79 208 -79 1 gnd
<< end >>
