magic
tech scmos
timestamp 1522765529
<< nwell >>
rect 5 113 184 139
rect 197 113 238 139
rect 253 113 294 139
rect 307 113 348 139
rect 101 8 188 34
rect 201 8 242 34
rect 257 8 298 34
rect 311 8 352 34
<< polysilicon >>
rect 42 126 44 128
rect 114 126 116 132
rect 153 126 155 132
rect 174 126 176 132
rect 207 126 209 132
rect 228 126 230 132
rect 263 126 265 132
rect 284 126 286 132
rect 317 126 319 132
rect 338 126 340 132
rect 42 109 44 120
rect 114 108 116 120
rect 153 108 155 120
rect 174 108 176 120
rect 207 108 209 120
rect 228 108 230 120
rect 263 108 265 120
rect 284 108 286 120
rect 317 108 319 120
rect 338 108 340 120
rect 42 87 44 105
rect 154 104 155 108
rect 175 104 176 108
rect 208 104 209 108
rect 229 104 230 108
rect 264 104 265 108
rect 285 104 286 108
rect 318 104 319 108
rect 339 104 340 108
rect 42 81 44 84
rect 114 86 116 104
rect 153 89 155 104
rect 174 89 176 104
rect 207 89 209 104
rect 228 89 230 104
rect 263 89 265 104
rect 284 89 286 104
rect 317 89 319 104
rect 338 89 340 104
rect 114 80 116 83
rect 153 80 155 83
rect 174 80 176 83
rect 207 80 209 83
rect 228 80 230 83
rect 263 80 265 83
rect 284 80 286 83
rect 317 80 319 83
rect 338 80 340 83
rect 118 64 120 67
rect 157 64 159 67
rect 178 64 180 67
rect 211 64 213 67
rect 232 64 234 67
rect 267 64 269 67
rect 288 64 290 67
rect 321 64 323 67
rect 342 64 344 67
rect 118 43 120 61
rect 157 43 159 58
rect 178 43 180 58
rect 211 43 213 58
rect 232 43 234 58
rect 267 43 269 58
rect 288 43 290 58
rect 321 43 323 58
rect 342 43 344 58
rect 158 39 159 43
rect 179 39 180 43
rect 212 39 213 43
rect 233 39 234 43
rect 268 39 269 43
rect 289 39 290 43
rect 322 39 323 43
rect 343 39 344 43
rect 118 27 120 39
rect 157 27 159 39
rect 178 27 180 39
rect 211 27 213 39
rect 232 27 234 39
rect 267 27 269 39
rect 288 27 290 39
rect 321 27 323 39
rect 342 27 344 39
rect 118 15 120 21
rect 157 15 159 21
rect 178 15 180 21
rect 211 15 213 21
rect 232 15 234 21
rect 267 15 269 21
rect 288 15 290 21
rect 321 15 323 21
rect 342 15 344 21
<< ndiffusion >>
rect 31 84 42 87
rect 44 84 61 87
rect 143 88 153 89
rect 103 83 114 86
rect 116 83 133 86
rect 143 84 145 88
rect 149 84 153 88
rect 143 83 153 84
rect 155 83 174 89
rect 176 88 184 89
rect 176 84 179 88
rect 183 84 184 88
rect 176 83 184 84
rect 197 88 207 89
rect 197 84 199 88
rect 203 84 207 88
rect 197 83 207 84
rect 209 83 228 89
rect 230 88 238 89
rect 230 84 233 88
rect 237 84 238 88
rect 230 83 238 84
rect 253 88 263 89
rect 253 84 255 88
rect 259 84 263 88
rect 253 83 263 84
rect 265 83 284 89
rect 286 88 294 89
rect 286 84 289 88
rect 293 84 294 88
rect 286 83 294 84
rect 307 88 317 89
rect 307 84 309 88
rect 313 84 317 88
rect 307 83 317 84
rect 319 83 338 89
rect 340 88 348 89
rect 340 84 343 88
rect 347 84 348 88
rect 340 83 348 84
rect 107 61 118 64
rect 120 61 137 64
rect 147 63 157 64
rect 147 59 149 63
rect 153 59 157 63
rect 147 58 157 59
rect 159 58 178 64
rect 180 63 188 64
rect 180 59 183 63
rect 187 59 188 63
rect 180 58 188 59
rect 201 63 211 64
rect 201 59 203 63
rect 207 59 211 63
rect 201 58 211 59
rect 213 58 232 64
rect 234 63 242 64
rect 234 59 237 63
rect 241 59 242 63
rect 234 58 242 59
rect 257 63 267 64
rect 257 59 259 63
rect 263 59 267 63
rect 257 58 267 59
rect 269 58 288 64
rect 290 63 298 64
rect 290 59 293 63
rect 297 59 298 63
rect 290 58 298 59
rect 311 63 321 64
rect 311 59 313 63
rect 317 59 321 63
rect 311 58 321 59
rect 323 58 342 64
rect 344 63 352 64
rect 344 59 347 63
rect 351 59 352 63
rect 344 58 352 59
<< pdiffusion >>
rect 11 125 42 126
rect 11 121 16 125
rect 20 121 42 125
rect 11 120 42 121
rect 44 121 60 126
rect 66 121 79 126
rect 44 120 79 121
rect 99 125 114 126
rect 103 121 114 125
rect 99 120 114 121
rect 116 125 136 126
rect 116 121 132 125
rect 116 120 136 121
rect 143 125 153 126
rect 143 121 145 125
rect 149 121 153 125
rect 143 120 153 121
rect 155 125 174 126
rect 155 121 162 125
rect 166 121 174 125
rect 155 120 174 121
rect 176 125 184 126
rect 176 121 179 125
rect 183 121 184 125
rect 176 120 184 121
rect 197 125 207 126
rect 197 121 199 125
rect 203 121 207 125
rect 197 120 207 121
rect 209 125 228 126
rect 209 121 216 125
rect 220 121 228 125
rect 209 120 228 121
rect 230 125 238 126
rect 230 121 233 125
rect 237 121 238 125
rect 230 120 238 121
rect 253 125 263 126
rect 253 121 255 125
rect 259 121 263 125
rect 253 120 263 121
rect 265 125 284 126
rect 265 121 272 125
rect 276 121 284 125
rect 265 120 284 121
rect 286 125 294 126
rect 286 121 289 125
rect 293 121 294 125
rect 286 120 294 121
rect 307 125 317 126
rect 307 121 309 125
rect 313 121 317 125
rect 307 120 317 121
rect 319 125 338 126
rect 319 121 326 125
rect 330 121 338 125
rect 319 120 338 121
rect 340 125 348 126
rect 340 121 343 125
rect 347 121 348 125
rect 340 120 348 121
rect 103 26 118 27
rect 107 22 118 26
rect 103 21 118 22
rect 120 26 140 27
rect 120 22 136 26
rect 120 21 140 22
rect 147 26 157 27
rect 147 22 149 26
rect 153 22 157 26
rect 147 21 157 22
rect 159 26 178 27
rect 159 22 166 26
rect 170 22 178 26
rect 159 21 178 22
rect 180 26 188 27
rect 180 22 183 26
rect 187 22 188 26
rect 180 21 188 22
rect 201 26 211 27
rect 201 22 203 26
rect 207 22 211 26
rect 201 21 211 22
rect 213 26 232 27
rect 213 22 220 26
rect 224 22 232 26
rect 213 21 232 22
rect 234 26 242 27
rect 234 22 237 26
rect 241 22 242 26
rect 234 21 242 22
rect 257 26 267 27
rect 257 22 259 26
rect 263 22 267 26
rect 257 21 267 22
rect 269 26 288 27
rect 269 22 276 26
rect 280 22 288 26
rect 269 21 288 22
rect 290 26 298 27
rect 290 22 293 26
rect 297 22 298 26
rect 290 21 298 22
rect 311 26 321 27
rect 311 22 313 26
rect 317 22 321 26
rect 311 21 321 22
rect 323 26 342 27
rect 323 22 330 26
rect 334 22 342 26
rect 323 21 342 22
rect 344 26 352 27
rect 344 22 347 26
rect 351 22 352 26
rect 344 21 352 22
<< metal1 >>
rect 0 144 366 147
rect 16 125 19 144
rect 61 127 65 129
rect 99 125 102 144
rect 162 125 165 144
rect 172 139 175 144
rect 216 125 219 144
rect 226 139 229 144
rect 272 125 275 144
rect 282 139 285 144
rect 326 125 329 144
rect 336 139 339 144
rect 61 110 65 121
rect 44 106 47 109
rect 61 100 64 110
rect 116 105 119 108
rect 61 96 62 100
rect 133 99 136 121
rect 146 116 149 121
rect 179 116 182 121
rect 146 113 182 116
rect 148 105 150 108
rect 170 105 171 108
rect 179 104 182 113
rect 200 116 203 121
rect 233 116 236 121
rect 200 113 236 116
rect 256 116 259 121
rect 289 116 292 121
rect 256 113 292 116
rect 310 116 313 121
rect 343 116 346 121
rect 310 113 346 116
rect 186 104 189 113
rect 200 108 207 109
rect 200 106 204 108
rect 221 104 225 107
rect 179 101 189 104
rect 61 88 64 96
rect 133 95 134 99
rect 133 87 136 95
rect 179 88 182 101
rect 221 100 224 104
rect 233 101 236 113
rect 289 112 292 113
rect 257 105 260 108
rect 233 98 252 101
rect 233 88 236 98
rect 281 102 284 104
rect 269 94 272 100
rect 283 98 284 102
rect 281 97 284 98
rect 246 91 272 94
rect 289 88 292 108
rect 313 104 314 107
rect 332 108 338 109
rect 332 106 335 108
rect 313 95 316 104
rect 343 103 346 113
rect 315 91 316 95
rect 343 88 346 99
rect 27 78 30 84
rect 99 78 102 83
rect 145 78 148 84
rect 199 78 202 84
rect 255 78 258 84
rect 309 78 312 84
rect 3 75 348 78
rect 171 72 176 75
rect 277 72 281 75
rect 103 69 352 72
rect 103 64 106 69
rect 149 63 152 69
rect 203 63 206 69
rect 259 63 262 69
rect 313 63 316 69
rect 137 52 140 60
rect 137 48 138 52
rect 120 39 123 42
rect 137 26 140 48
rect 183 46 186 59
rect 183 43 193 46
rect 225 43 228 47
rect 237 49 240 59
rect 237 46 256 49
rect 285 49 288 50
rect 152 39 154 42
rect 174 39 175 42
rect 183 34 186 43
rect 150 31 186 34
rect 150 26 153 31
rect 183 26 186 31
rect 190 34 193 43
rect 204 39 208 41
rect 225 40 229 43
rect 204 38 211 39
rect 237 34 240 46
rect 287 45 288 49
rect 285 43 288 45
rect 261 39 264 42
rect 293 39 296 59
rect 319 52 320 56
rect 317 43 320 52
rect 347 48 350 59
rect 317 40 318 43
rect 336 39 339 41
rect 336 38 342 39
rect 293 34 296 35
rect 347 34 350 44
rect 204 31 240 34
rect 204 26 207 31
rect 237 26 240 31
rect 260 31 296 34
rect 260 26 263 31
rect 293 26 296 31
rect 314 31 350 34
rect 314 26 317 31
rect 347 26 350 31
rect 103 3 106 22
rect 166 3 169 22
rect 176 3 179 8
rect 220 3 223 22
rect 230 3 233 8
rect 276 3 279 22
rect 286 3 289 8
rect 330 3 333 22
rect 340 3 343 8
rect 361 3 366 144
rect 101 0 366 3
<< metal2 >>
rect 90 116 170 119
rect 90 110 93 116
rect 51 107 93 110
rect 166 109 169 116
rect 190 114 249 117
rect 123 106 144 109
rect 170 106 196 109
rect 200 106 201 109
rect 246 108 249 114
rect 270 109 289 112
rect 246 105 253 108
rect 270 104 273 109
rect 293 110 332 111
rect 293 108 328 110
rect 66 96 78 99
rect 75 32 78 96
rect 138 96 220 99
rect 283 99 342 102
rect 253 94 256 97
rect 253 91 311 94
rect 242 72 246 90
rect 123 68 246 72
rect 123 42 127 68
rect 242 67 246 68
rect 257 53 315 56
rect 142 48 224 51
rect 257 50 260 53
rect 287 45 346 48
rect 127 38 148 41
rect 174 38 200 41
rect 204 38 205 41
rect 250 39 257 42
rect 170 32 173 38
rect 75 29 173 32
rect 250 33 253 39
rect 297 37 332 39
rect 297 36 336 37
rect 194 30 253 33
<< ntransistor >>
rect 42 84 44 87
rect 114 83 116 86
rect 153 83 155 89
rect 174 83 176 89
rect 207 83 209 89
rect 228 83 230 89
rect 263 83 265 89
rect 284 83 286 89
rect 317 83 319 89
rect 338 83 340 89
rect 118 61 120 64
rect 157 58 159 64
rect 178 58 180 64
rect 211 58 213 64
rect 232 58 234 64
rect 267 58 269 64
rect 288 58 290 64
rect 321 58 323 64
rect 342 58 344 64
<< ptransistor >>
rect 42 120 44 126
rect 114 120 116 126
rect 153 120 155 126
rect 174 120 176 126
rect 207 120 209 126
rect 228 120 230 126
rect 263 120 265 126
rect 284 120 286 126
rect 317 120 319 126
rect 338 120 340 126
rect 118 21 120 27
rect 157 21 159 27
rect 178 21 180 27
rect 211 21 213 27
rect 232 21 234 27
rect 267 21 269 27
rect 288 21 290 27
rect 321 21 323 27
rect 342 21 344 27
<< polycontact >>
rect 40 105 44 109
rect 112 104 116 108
rect 150 104 154 108
rect 171 104 175 108
rect 204 104 208 108
rect 225 104 229 108
rect 260 104 264 108
rect 281 104 285 108
rect 314 104 318 108
rect 335 104 339 108
rect 116 39 120 43
rect 154 39 158 43
rect 175 39 179 43
rect 208 39 212 43
rect 229 39 233 43
rect 264 39 268 43
rect 285 39 289 43
rect 318 39 322 43
rect 339 39 343 43
<< ndcontact >>
rect 27 84 31 88
rect 61 84 65 88
rect 99 83 103 87
rect 133 83 137 87
rect 145 84 149 88
rect 179 84 183 88
rect 199 84 203 88
rect 233 84 237 88
rect 255 84 259 88
rect 289 84 293 88
rect 309 84 313 88
rect 343 84 347 88
rect 103 60 107 64
rect 137 60 141 64
rect 149 59 153 63
rect 183 59 187 63
rect 203 59 207 63
rect 237 59 241 63
rect 259 59 263 63
rect 293 59 297 63
rect 313 59 317 63
rect 347 59 351 63
<< pdcontact >>
rect 16 121 20 125
rect 60 121 66 127
rect 99 121 103 125
rect 132 121 136 125
rect 145 121 149 125
rect 162 121 166 125
rect 179 121 183 125
rect 199 121 203 125
rect 216 121 220 125
rect 233 121 237 125
rect 255 121 259 125
rect 272 121 276 125
rect 289 121 293 125
rect 309 121 313 125
rect 326 121 330 125
rect 343 121 347 125
rect 103 22 107 26
rect 136 22 140 26
rect 149 22 153 26
rect 166 22 170 26
rect 183 22 187 26
rect 203 22 207 26
rect 220 22 224 26
rect 237 22 241 26
rect 259 22 263 26
rect 276 22 280 26
rect 293 22 297 26
rect 313 22 317 26
rect 330 22 334 26
rect 347 22 351 26
<< m2contact >>
rect 47 106 51 110
rect 119 105 123 109
rect 62 96 66 100
rect 144 105 148 109
rect 166 105 170 109
rect 186 113 190 117
rect 196 105 200 109
rect 134 95 138 99
rect 220 96 224 100
rect 253 105 257 109
rect 289 108 293 112
rect 252 97 256 101
rect 269 100 273 104
rect 279 98 283 102
rect 242 90 246 94
rect 328 106 332 110
rect 342 99 346 103
rect 311 91 315 95
rect 138 48 142 52
rect 123 38 127 42
rect 224 47 228 51
rect 256 46 260 50
rect 148 38 152 42
rect 170 38 174 42
rect 200 38 204 42
rect 283 45 287 49
rect 257 38 261 42
rect 315 52 319 56
rect 346 44 350 48
rect 293 35 297 39
rect 332 37 336 41
rect 190 30 194 34
<< nsubstratencontact >>
rect 172 135 176 139
rect 226 135 230 139
rect 282 135 286 139
rect 336 135 340 139
rect 176 8 180 12
rect 230 8 234 12
rect 286 8 290 12
rect 340 8 344 12
<< labels >>
rlabel metal1 328 76 328 76 1 gnd
rlabel metal1 332 2 332 2 1 vdd
rlabel metal1 332 71 332 71 5 gnd
rlabel m2contact 63 98 63 98 1 en_bar_D2
rlabel polycontact 152 106 152 106 1 D_D2
rlabel metal1 134 105 134 105 1 D_bar_D2
rlabel ndiffusion 162 86 162 86 1 n1_D2
rlabel polycontact 173 106 173 106 1 en_D2
rlabel metal1 181 103 181 103 1 out_n1_D2
rlabel ndiffusion 218 86 218 86 1 n2_D2
rlabel metal1 236 99 236 99 1 out_n2_D2
rlabel ndiffusion 274 86 274 86 1 n3_D2
rlabel ndiffusion 328 86 328 86 1 n4_D2
rlabel m2contact 349 45 349 45 1 q_bar_D2
rlabel ndiffusion 332 61 332 61 1 n10_D2
rlabel m2contact 295 37 295 37 1 q_D2
rlabel ndiffusion 278 61 278 61 1 n9_D2
rlabel metal1 240 48 240 48 1 out_n8_D2
rlabel ndiffusion 222 61 222 61 1 n8_D2
rlabel metal1 185 44 185 44 1 out_n7__D2
rlabel ndiffusion 166 61 166 61 1 n7_D2
rlabel polycontact 156 41 156 41 1 q_l1_D2
rlabel metal1 138 45 138 45 1 n6_D2
rlabel m2contact 345 102 345 102 1 q_l1_bar_D2
<< end >>
