magic
tech scmos
timestamp 1523034434
<< nwell >>
rect 37 80 216 106
rect 229 80 270 106
rect 285 80 326 106
rect 339 80 380 106
rect 133 -25 220 1
rect 233 -25 274 1
rect 289 -25 330 1
rect 343 -25 384 1
<< polysilicon >>
rect 74 93 76 95
rect 146 93 148 99
rect 185 93 187 99
rect 206 93 208 99
rect 239 93 241 99
rect 260 93 262 99
rect 295 93 297 99
rect 316 93 318 99
rect 349 93 351 99
rect 370 93 372 99
rect 74 76 76 87
rect 146 75 148 87
rect 185 75 187 87
rect 206 75 208 87
rect 239 75 241 87
rect 260 75 262 87
rect 295 75 297 87
rect 316 75 318 87
rect 349 75 351 87
rect 370 75 372 87
rect 74 54 76 72
rect 186 71 187 75
rect 207 71 208 75
rect 240 71 241 75
rect 261 71 262 75
rect 296 71 297 75
rect 317 71 318 75
rect 350 71 351 75
rect 371 71 372 75
rect 74 48 76 51
rect 146 53 148 71
rect 185 56 187 71
rect 206 56 208 71
rect 239 56 241 71
rect 260 56 262 71
rect 295 56 297 71
rect 316 56 318 71
rect 349 56 351 71
rect 370 56 372 71
rect 146 47 148 50
rect 185 47 187 50
rect 206 47 208 50
rect 239 47 241 50
rect 260 47 262 50
rect 295 47 297 50
rect 316 47 318 50
rect 349 47 351 50
rect 370 47 372 50
rect 150 31 152 34
rect 189 31 191 34
rect 210 31 212 34
rect 243 31 245 34
rect 264 31 266 34
rect 299 31 301 34
rect 320 31 322 34
rect 353 31 355 34
rect 374 31 376 34
rect 150 10 152 28
rect 189 10 191 25
rect 210 10 212 25
rect 243 10 245 25
rect 264 10 266 25
rect 299 10 301 25
rect 320 10 322 25
rect 353 10 355 25
rect 374 10 376 25
rect 190 6 191 10
rect 211 6 212 10
rect 244 6 245 10
rect 265 6 266 10
rect 300 6 301 10
rect 321 6 322 10
rect 354 6 355 10
rect 375 6 376 10
rect 150 -6 152 6
rect 189 -6 191 6
rect 210 -6 212 6
rect 243 -6 245 6
rect 264 -6 266 6
rect 299 -6 301 6
rect 320 -6 322 6
rect 353 -6 355 6
rect 374 -6 376 6
rect 150 -18 152 -12
rect 189 -18 191 -12
rect 210 -18 212 -12
rect 243 -18 245 -12
rect 264 -18 266 -12
rect 299 -18 301 -12
rect 320 -18 322 -12
rect 353 -18 355 -12
rect 374 -18 376 -12
<< ndiffusion >>
rect 63 51 74 54
rect 76 51 93 54
rect 175 55 185 56
rect 135 50 146 53
rect 148 50 165 53
rect 175 51 177 55
rect 181 51 185 55
rect 175 50 185 51
rect 187 50 206 56
rect 208 55 216 56
rect 208 51 211 55
rect 215 51 216 55
rect 208 50 216 51
rect 229 55 239 56
rect 229 51 231 55
rect 235 51 239 55
rect 229 50 239 51
rect 241 50 260 56
rect 262 55 270 56
rect 262 51 265 55
rect 269 51 270 55
rect 262 50 270 51
rect 285 55 295 56
rect 285 51 287 55
rect 291 51 295 55
rect 285 50 295 51
rect 297 50 316 56
rect 318 55 326 56
rect 318 51 321 55
rect 325 51 326 55
rect 318 50 326 51
rect 339 55 349 56
rect 339 51 341 55
rect 345 51 349 55
rect 339 50 349 51
rect 351 50 370 56
rect 372 55 380 56
rect 372 51 375 55
rect 379 51 380 55
rect 372 50 380 51
rect 139 28 150 31
rect 152 28 169 31
rect 179 30 189 31
rect 179 26 181 30
rect 185 26 189 30
rect 179 25 189 26
rect 191 25 210 31
rect 212 30 220 31
rect 212 26 215 30
rect 219 26 220 30
rect 212 25 220 26
rect 233 30 243 31
rect 233 26 235 30
rect 239 26 243 30
rect 233 25 243 26
rect 245 25 264 31
rect 266 30 274 31
rect 266 26 269 30
rect 273 26 274 30
rect 266 25 274 26
rect 289 30 299 31
rect 289 26 291 30
rect 295 26 299 30
rect 289 25 299 26
rect 301 25 320 31
rect 322 30 330 31
rect 322 26 325 30
rect 329 26 330 30
rect 322 25 330 26
rect 343 30 353 31
rect 343 26 345 30
rect 349 26 353 30
rect 343 25 353 26
rect 355 25 374 31
rect 376 30 384 31
rect 376 26 379 30
rect 383 26 384 30
rect 376 25 384 26
<< pdiffusion >>
rect 43 92 74 93
rect 43 88 48 92
rect 52 88 74 92
rect 43 87 74 88
rect 76 88 92 93
rect 98 88 111 93
rect 76 87 111 88
rect 131 92 146 93
rect 135 88 146 92
rect 131 87 146 88
rect 148 92 168 93
rect 148 88 164 92
rect 148 87 168 88
rect 175 92 185 93
rect 175 88 177 92
rect 181 88 185 92
rect 175 87 185 88
rect 187 92 206 93
rect 187 88 194 92
rect 198 88 206 92
rect 187 87 206 88
rect 208 92 216 93
rect 208 88 211 92
rect 215 88 216 92
rect 208 87 216 88
rect 229 92 239 93
rect 229 88 231 92
rect 235 88 239 92
rect 229 87 239 88
rect 241 92 260 93
rect 241 88 248 92
rect 252 88 260 92
rect 241 87 260 88
rect 262 92 270 93
rect 262 88 265 92
rect 269 88 270 92
rect 262 87 270 88
rect 285 92 295 93
rect 285 88 287 92
rect 291 88 295 92
rect 285 87 295 88
rect 297 92 316 93
rect 297 88 304 92
rect 308 88 316 92
rect 297 87 316 88
rect 318 92 326 93
rect 318 88 321 92
rect 325 88 326 92
rect 318 87 326 88
rect 339 92 349 93
rect 339 88 341 92
rect 345 88 349 92
rect 339 87 349 88
rect 351 92 370 93
rect 351 88 358 92
rect 362 88 370 92
rect 351 87 370 88
rect 372 92 380 93
rect 372 88 375 92
rect 379 88 380 92
rect 372 87 380 88
rect 135 -7 150 -6
rect 139 -11 150 -7
rect 135 -12 150 -11
rect 152 -7 172 -6
rect 152 -11 168 -7
rect 152 -12 172 -11
rect 179 -7 189 -6
rect 179 -11 181 -7
rect 185 -11 189 -7
rect 179 -12 189 -11
rect 191 -7 210 -6
rect 191 -11 198 -7
rect 202 -11 210 -7
rect 191 -12 210 -11
rect 212 -7 220 -6
rect 212 -11 215 -7
rect 219 -11 220 -7
rect 212 -12 220 -11
rect 233 -7 243 -6
rect 233 -11 235 -7
rect 239 -11 243 -7
rect 233 -12 243 -11
rect 245 -7 264 -6
rect 245 -11 252 -7
rect 256 -11 264 -7
rect 245 -12 264 -11
rect 266 -7 274 -6
rect 266 -11 269 -7
rect 273 -11 274 -7
rect 266 -12 274 -11
rect 289 -7 299 -6
rect 289 -11 291 -7
rect 295 -11 299 -7
rect 289 -12 299 -11
rect 301 -7 320 -6
rect 301 -11 308 -7
rect 312 -11 320 -7
rect 301 -12 320 -11
rect 322 -7 330 -6
rect 322 -11 325 -7
rect 329 -11 330 -7
rect 322 -12 330 -11
rect 343 -7 353 -6
rect 343 -11 345 -7
rect 349 -11 353 -7
rect 343 -12 353 -11
rect 355 -7 374 -6
rect 355 -11 362 -7
rect 366 -11 374 -7
rect 355 -12 374 -11
rect 376 -7 384 -6
rect 376 -11 379 -7
rect 383 -11 384 -7
rect 376 -12 384 -11
<< metal1 >>
rect 32 111 398 114
rect 48 92 51 111
rect 93 94 97 96
rect 131 92 134 111
rect 194 92 197 111
rect 204 106 207 111
rect 248 92 251 111
rect 258 106 261 111
rect 304 92 307 111
rect 314 106 317 111
rect 358 92 361 111
rect 368 106 371 111
rect 93 77 97 88
rect 76 73 79 76
rect 93 67 96 77
rect 148 72 151 75
rect 93 63 94 67
rect 165 66 168 88
rect 178 83 181 88
rect 211 83 214 88
rect 178 80 214 83
rect 180 72 182 75
rect 202 72 203 75
rect 211 71 214 80
rect 232 83 235 88
rect 265 83 268 88
rect 232 80 268 83
rect 288 83 291 88
rect 321 83 324 88
rect 288 80 324 83
rect 342 83 345 88
rect 375 83 378 88
rect 342 80 378 83
rect 218 71 221 80
rect 232 75 239 76
rect 232 73 236 75
rect 253 71 257 74
rect 211 68 221 71
rect 93 55 96 63
rect 165 62 166 66
rect 165 54 168 62
rect 211 55 214 68
rect 253 67 256 71
rect 265 68 268 80
rect 321 79 324 80
rect 289 72 292 75
rect 265 65 284 68
rect 265 55 268 65
rect 313 69 316 71
rect 301 61 304 67
rect 315 65 316 69
rect 313 64 316 65
rect 278 58 304 61
rect 321 55 324 75
rect 345 71 346 74
rect 364 75 370 76
rect 364 73 367 75
rect 345 62 348 71
rect 375 70 378 80
rect 347 58 348 62
rect 375 55 378 66
rect 59 45 62 51
rect 131 45 134 50
rect 177 45 180 51
rect 231 45 234 51
rect 287 45 290 51
rect 341 45 344 51
rect 35 42 380 45
rect 203 39 208 42
rect 309 39 313 42
rect 135 36 384 39
rect 135 31 138 36
rect 181 30 184 36
rect 235 30 238 36
rect 291 30 294 36
rect 345 30 348 36
rect 169 19 172 27
rect 169 15 170 19
rect 152 6 155 9
rect 169 -7 172 15
rect 215 13 218 26
rect 215 10 225 13
rect 257 10 260 14
rect 269 16 272 26
rect 269 13 288 16
rect 317 16 320 17
rect 184 6 186 9
rect 206 6 207 9
rect 215 1 218 10
rect 182 -2 218 1
rect 182 -7 185 -2
rect 215 -7 218 -2
rect 222 1 225 10
rect 236 6 240 8
rect 257 7 261 10
rect 236 5 243 6
rect 269 1 272 13
rect 319 12 320 16
rect 317 10 320 12
rect 293 6 296 9
rect 325 6 328 26
rect 351 19 352 23
rect 349 10 352 19
rect 379 15 382 26
rect 349 7 350 10
rect 368 6 371 8
rect 368 5 374 6
rect 325 1 328 2
rect 379 1 382 11
rect 236 -2 272 1
rect 236 -7 239 -2
rect 269 -7 272 -2
rect 292 -2 328 1
rect 292 -7 295 -2
rect 325 -7 328 -2
rect 346 -2 382 1
rect 346 -7 349 -2
rect 379 -7 382 -2
rect 135 -30 138 -11
rect 198 -30 201 -11
rect 208 -30 211 -25
rect 252 -30 255 -11
rect 262 -30 265 -25
rect 308 -30 311 -11
rect 318 -30 321 -25
rect 362 -30 365 -11
rect 372 -30 375 -25
rect 393 -30 398 111
rect 133 -33 398 -30
<< metal2 >>
rect 122 83 202 86
rect 122 77 125 83
rect 83 74 125 77
rect 198 76 201 83
rect 222 81 281 84
rect 155 73 176 76
rect 202 73 228 76
rect 232 73 233 76
rect 278 75 281 81
rect 302 76 321 79
rect 278 72 285 75
rect 302 71 305 76
rect 325 77 364 78
rect 325 75 360 77
rect 98 63 110 66
rect 107 -1 110 63
rect 170 63 252 66
rect 315 66 374 69
rect 285 61 288 64
rect 285 58 343 61
rect 274 39 278 57
rect 155 35 278 39
rect 155 9 159 35
rect 274 34 278 35
rect 289 20 347 23
rect 174 15 256 18
rect 289 17 292 20
rect 319 12 378 15
rect 159 5 180 8
rect 206 5 232 8
rect 236 5 237 8
rect 282 6 289 9
rect 202 -1 205 5
rect 107 -4 205 -1
rect 282 0 285 6
rect 329 4 364 6
rect 329 3 368 4
rect 226 -3 285 0
<< ntransistor >>
rect 74 51 76 54
rect 146 50 148 53
rect 185 50 187 56
rect 206 50 208 56
rect 239 50 241 56
rect 260 50 262 56
rect 295 50 297 56
rect 316 50 318 56
rect 349 50 351 56
rect 370 50 372 56
rect 150 28 152 31
rect 189 25 191 31
rect 210 25 212 31
rect 243 25 245 31
rect 264 25 266 31
rect 299 25 301 31
rect 320 25 322 31
rect 353 25 355 31
rect 374 25 376 31
<< ptransistor >>
rect 74 87 76 93
rect 146 87 148 93
rect 185 87 187 93
rect 206 87 208 93
rect 239 87 241 93
rect 260 87 262 93
rect 295 87 297 93
rect 316 87 318 93
rect 349 87 351 93
rect 370 87 372 93
rect 150 -12 152 -6
rect 189 -12 191 -6
rect 210 -12 212 -6
rect 243 -12 245 -6
rect 264 -12 266 -6
rect 299 -12 301 -6
rect 320 -12 322 -6
rect 353 -12 355 -6
rect 374 -12 376 -6
<< polycontact >>
rect 72 72 76 76
rect 144 71 148 75
rect 182 71 186 75
rect 203 71 207 75
rect 236 71 240 75
rect 257 71 261 75
rect 292 71 296 75
rect 313 71 317 75
rect 346 71 350 75
rect 367 71 371 75
rect 148 6 152 10
rect 186 6 190 10
rect 207 6 211 10
rect 240 6 244 10
rect 261 6 265 10
rect 296 6 300 10
rect 317 6 321 10
rect 350 6 354 10
rect 371 6 375 10
<< ndcontact >>
rect 59 51 63 55
rect 93 51 97 55
rect 131 50 135 54
rect 165 50 169 54
rect 177 51 181 55
rect 211 51 215 55
rect 231 51 235 55
rect 265 51 269 55
rect 287 51 291 55
rect 321 51 325 55
rect 341 51 345 55
rect 375 51 379 55
rect 135 27 139 31
rect 169 27 173 31
rect 181 26 185 30
rect 215 26 219 30
rect 235 26 239 30
rect 269 26 273 30
rect 291 26 295 30
rect 325 26 329 30
rect 345 26 349 30
rect 379 26 383 30
<< pdcontact >>
rect 48 88 52 92
rect 92 88 98 94
rect 131 88 135 92
rect 164 88 168 92
rect 177 88 181 92
rect 194 88 198 92
rect 211 88 215 92
rect 231 88 235 92
rect 248 88 252 92
rect 265 88 269 92
rect 287 88 291 92
rect 304 88 308 92
rect 321 88 325 92
rect 341 88 345 92
rect 358 88 362 92
rect 375 88 379 92
rect 135 -11 139 -7
rect 168 -11 172 -7
rect 181 -11 185 -7
rect 198 -11 202 -7
rect 215 -11 219 -7
rect 235 -11 239 -7
rect 252 -11 256 -7
rect 269 -11 273 -7
rect 291 -11 295 -7
rect 308 -11 312 -7
rect 325 -11 329 -7
rect 345 -11 349 -7
rect 362 -11 366 -7
rect 379 -11 383 -7
<< m2contact >>
rect 79 73 83 77
rect 151 72 155 76
rect 94 63 98 67
rect 176 72 180 76
rect 198 72 202 76
rect 218 80 222 84
rect 228 72 232 76
rect 166 62 170 66
rect 252 63 256 67
rect 285 72 289 76
rect 321 75 325 79
rect 284 64 288 68
rect 301 67 305 71
rect 311 65 315 69
rect 274 57 278 61
rect 360 73 364 77
rect 374 66 378 70
rect 343 58 347 62
rect 170 15 174 19
rect 155 5 159 9
rect 256 14 260 18
rect 288 13 292 17
rect 180 5 184 9
rect 202 5 206 9
rect 232 5 236 9
rect 315 12 319 16
rect 289 5 293 9
rect 347 19 351 23
rect 378 11 382 15
rect 325 2 329 6
rect 364 4 368 8
rect 222 -3 226 1
<< nsubstratencontact >>
rect 204 102 208 106
rect 258 102 262 106
rect 314 102 318 106
rect 368 102 372 106
rect 208 -25 212 -21
rect 262 -25 266 -21
rect 318 -25 322 -21
rect 372 -25 376 -21
<< labels >>
rlabel metal1 364 -31 364 -31 1 vdd
rlabel m2contact 95 65 95 65 1 en_bar_D4
rlabel metal1 166 72 166 72 1 D_bar_D4
rlabel polycontact 184 73 184 73 1 D_D4
rlabel polycontact 205 73 205 73 1 en_D4
rlabel ndiffusion 194 53 194 53 1 n1_D4
rlabel ndiffusion 250 53 250 53 1 n2_D4
rlabel metal1 268 66 268 66 1 out_n2_D4
rlabel ndiffusion 306 53 306 53 1 n3_D4
rlabel ndiffusion 360 53 360 53 1 n4_D4
rlabel m2contact 375 68 375 68 1 q_l1_bar_D4
rlabel metal1 311 42 311 42 1 vss
rlabel ndiffusion 364 28 364 28 1 n10_D4
rlabel m2contact 381 12 381 12 1 q_bar_D4
rlabel m2contact 327 4 327 4 1 q_D4
rlabel ndiffusion 310 28 310 28 1 n9_D4
rlabel ndiffusion 254 28 254 28 1 n8_D4
rlabel metal1 272 15 272 15 1 out_n8_D4
rlabel metal1 217 11 217 11 1 out_n7_D4
rlabel ndiffusion 198 28 198 28 1 n7_D4
rlabel polycontact 188 8 188 8 1 q_l1_D4
rlabel metal1 170 12 170 12 1 n6_D4
rlabel metal1 213 70 213 70 1 out_n1_D4
<< end >>
