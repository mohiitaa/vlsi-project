magic
tech scmos
timestamp 1522727561
<< nwell >>
rect -92 38 87 64
rect 100 38 141 64
rect 156 38 197 64
rect 210 38 251 64
rect 4 -67 91 -41
rect 104 -67 145 -41
rect 160 -67 201 -41
rect 214 -67 255 -41
<< polysilicon >>
rect -55 51 -53 53
rect 17 51 19 57
rect 56 51 58 57
rect 77 51 79 57
rect 110 51 112 57
rect 131 51 133 57
rect 166 51 168 57
rect 187 51 189 57
rect 220 51 222 57
rect 241 51 243 57
rect -55 34 -53 45
rect 17 33 19 45
rect 56 33 58 45
rect 77 33 79 45
rect 110 33 112 45
rect 131 33 133 45
rect 166 33 168 45
rect 187 33 189 45
rect 220 33 222 45
rect 241 33 243 45
rect -55 12 -53 30
rect 57 29 58 33
rect 78 29 79 33
rect 111 29 112 33
rect 132 29 133 33
rect 167 29 168 33
rect 188 29 189 33
rect 221 29 222 33
rect 242 29 243 33
rect -55 6 -53 9
rect 17 11 19 29
rect 56 14 58 29
rect 77 14 79 29
rect 110 14 112 29
rect 131 14 133 29
rect 166 14 168 29
rect 187 14 189 29
rect 220 14 222 29
rect 241 14 243 29
rect 17 5 19 8
rect 56 5 58 8
rect 77 5 79 8
rect 110 5 112 8
rect 131 5 133 8
rect 166 5 168 8
rect 187 5 189 8
rect 220 5 222 8
rect 241 5 243 8
rect 21 -11 23 -8
rect 60 -11 62 -8
rect 81 -11 83 -8
rect 114 -11 116 -8
rect 135 -11 137 -8
rect 170 -11 172 -8
rect 191 -11 193 -8
rect 224 -11 226 -8
rect 245 -11 247 -8
rect 21 -32 23 -14
rect 60 -32 62 -17
rect 81 -32 83 -17
rect 114 -32 116 -17
rect 135 -32 137 -17
rect 170 -32 172 -17
rect 191 -32 193 -17
rect 224 -32 226 -17
rect 245 -32 247 -17
rect 61 -36 62 -32
rect 82 -36 83 -32
rect 115 -36 116 -32
rect 136 -36 137 -32
rect 171 -36 172 -32
rect 192 -36 193 -32
rect 225 -36 226 -32
rect 246 -36 247 -32
rect 21 -48 23 -36
rect 60 -48 62 -36
rect 81 -48 83 -36
rect 114 -48 116 -36
rect 135 -48 137 -36
rect 170 -48 172 -36
rect 191 -48 193 -36
rect 224 -48 226 -36
rect 245 -48 247 -36
rect 21 -60 23 -54
rect 60 -60 62 -54
rect 81 -60 83 -54
rect 114 -60 116 -54
rect 135 -60 137 -54
rect 170 -60 172 -54
rect 191 -60 193 -54
rect 224 -60 226 -54
rect 245 -60 247 -54
<< ndiffusion >>
rect -66 9 -55 12
rect -53 9 -36 12
rect 46 13 56 14
rect 6 8 17 11
rect 19 8 36 11
rect 46 9 48 13
rect 52 9 56 13
rect 46 8 56 9
rect 58 8 77 14
rect 79 13 87 14
rect 79 9 82 13
rect 86 9 87 13
rect 79 8 87 9
rect 100 13 110 14
rect 100 9 102 13
rect 106 9 110 13
rect 100 8 110 9
rect 112 8 131 14
rect 133 13 141 14
rect 133 9 136 13
rect 140 9 141 13
rect 133 8 141 9
rect 156 13 166 14
rect 156 9 158 13
rect 162 9 166 13
rect 156 8 166 9
rect 168 8 187 14
rect 189 13 197 14
rect 189 9 192 13
rect 196 9 197 13
rect 189 8 197 9
rect 210 13 220 14
rect 210 9 212 13
rect 216 9 220 13
rect 210 8 220 9
rect 222 8 241 14
rect 243 13 251 14
rect 243 9 246 13
rect 250 9 251 13
rect 243 8 251 9
rect 10 -14 21 -11
rect 23 -14 40 -11
rect 50 -12 60 -11
rect 50 -16 52 -12
rect 56 -16 60 -12
rect 50 -17 60 -16
rect 62 -17 81 -11
rect 83 -12 91 -11
rect 83 -16 86 -12
rect 90 -16 91 -12
rect 83 -17 91 -16
rect 104 -12 114 -11
rect 104 -16 106 -12
rect 110 -16 114 -12
rect 104 -17 114 -16
rect 116 -17 135 -11
rect 137 -12 145 -11
rect 137 -16 140 -12
rect 144 -16 145 -12
rect 137 -17 145 -16
rect 160 -12 170 -11
rect 160 -16 162 -12
rect 166 -16 170 -12
rect 160 -17 170 -16
rect 172 -17 191 -11
rect 193 -12 201 -11
rect 193 -16 196 -12
rect 200 -16 201 -12
rect 193 -17 201 -16
rect 214 -12 224 -11
rect 214 -16 216 -12
rect 220 -16 224 -12
rect 214 -17 224 -16
rect 226 -17 245 -11
rect 247 -12 255 -11
rect 247 -16 250 -12
rect 254 -16 255 -12
rect 247 -17 255 -16
<< pdiffusion >>
rect -86 50 -55 51
rect -86 46 -81 50
rect -77 46 -55 50
rect -86 45 -55 46
rect -53 46 -37 51
rect -31 46 -18 51
rect -53 45 -18 46
rect 2 50 17 51
rect 6 46 17 50
rect 2 45 17 46
rect 19 50 39 51
rect 19 46 35 50
rect 19 45 39 46
rect 46 50 56 51
rect 46 46 48 50
rect 52 46 56 50
rect 46 45 56 46
rect 58 50 77 51
rect 58 46 65 50
rect 69 46 77 50
rect 58 45 77 46
rect 79 50 87 51
rect 79 46 82 50
rect 86 46 87 50
rect 79 45 87 46
rect 100 50 110 51
rect 100 46 102 50
rect 106 46 110 50
rect 100 45 110 46
rect 112 50 131 51
rect 112 46 119 50
rect 123 46 131 50
rect 112 45 131 46
rect 133 50 141 51
rect 133 46 136 50
rect 140 46 141 50
rect 133 45 141 46
rect 156 50 166 51
rect 156 46 158 50
rect 162 46 166 50
rect 156 45 166 46
rect 168 50 187 51
rect 168 46 175 50
rect 179 46 187 50
rect 168 45 187 46
rect 189 50 197 51
rect 189 46 192 50
rect 196 46 197 50
rect 189 45 197 46
rect 210 50 220 51
rect 210 46 212 50
rect 216 46 220 50
rect 210 45 220 46
rect 222 50 241 51
rect 222 46 229 50
rect 233 46 241 50
rect 222 45 241 46
rect 243 50 251 51
rect 243 46 246 50
rect 250 46 251 50
rect 243 45 251 46
rect 6 -49 21 -48
rect 10 -53 21 -49
rect 6 -54 21 -53
rect 23 -49 43 -48
rect 23 -53 39 -49
rect 23 -54 43 -53
rect 50 -49 60 -48
rect 50 -53 52 -49
rect 56 -53 60 -49
rect 50 -54 60 -53
rect 62 -49 81 -48
rect 62 -53 69 -49
rect 73 -53 81 -49
rect 62 -54 81 -53
rect 83 -49 91 -48
rect 83 -53 86 -49
rect 90 -53 91 -49
rect 83 -54 91 -53
rect 104 -49 114 -48
rect 104 -53 106 -49
rect 110 -53 114 -49
rect 104 -54 114 -53
rect 116 -49 135 -48
rect 116 -53 123 -49
rect 127 -53 135 -49
rect 116 -54 135 -53
rect 137 -49 145 -48
rect 137 -53 140 -49
rect 144 -53 145 -49
rect 137 -54 145 -53
rect 160 -49 170 -48
rect 160 -53 162 -49
rect 166 -53 170 -49
rect 160 -54 170 -53
rect 172 -49 191 -48
rect 172 -53 179 -49
rect 183 -53 191 -49
rect 172 -54 191 -53
rect 193 -49 201 -48
rect 193 -53 196 -49
rect 200 -53 201 -49
rect 193 -54 201 -53
rect 214 -49 224 -48
rect 214 -53 216 -49
rect 220 -53 224 -49
rect 214 -54 224 -53
rect 226 -49 245 -48
rect 226 -53 233 -49
rect 237 -53 245 -49
rect 226 -54 245 -53
rect 247 -49 255 -48
rect 247 -53 250 -49
rect 254 -53 255 -49
rect 247 -54 255 -53
<< metal1 >>
rect -97 69 269 72
rect -81 50 -78 69
rect -36 52 -32 54
rect 2 50 5 69
rect 65 50 68 69
rect 75 64 78 69
rect 119 50 122 69
rect 129 64 132 69
rect 175 50 178 69
rect 185 64 188 69
rect 229 50 232 69
rect 239 64 242 69
rect -36 35 -32 46
rect -53 31 -50 34
rect -36 25 -33 35
rect 19 30 22 33
rect -36 21 -35 25
rect 36 24 39 46
rect 49 41 52 46
rect 82 41 85 46
rect 49 38 85 41
rect 51 30 53 33
rect 73 30 74 33
rect 82 29 85 38
rect 103 41 106 46
rect 136 41 139 46
rect 103 38 139 41
rect 159 41 162 46
rect 192 41 195 46
rect 159 38 195 41
rect 213 41 216 46
rect 246 41 249 46
rect 213 38 249 41
rect 89 29 92 38
rect 103 33 110 34
rect 103 31 107 33
rect 124 29 128 32
rect 82 26 92 29
rect -36 13 -33 21
rect 36 20 37 24
rect 36 12 39 20
rect 82 13 85 26
rect 124 25 127 29
rect 136 26 139 38
rect 192 37 195 38
rect 160 30 163 33
rect 136 23 155 26
rect 136 13 139 23
rect 184 27 187 29
rect 172 19 175 25
rect 186 23 187 27
rect 184 22 187 23
rect 149 16 175 19
rect 192 13 195 33
rect 216 29 217 32
rect 235 33 241 34
rect 235 31 238 33
rect 216 20 219 29
rect 246 28 249 38
rect 218 16 219 20
rect 246 13 249 24
rect -70 3 -67 9
rect 2 3 5 8
rect 48 3 51 9
rect 102 3 105 9
rect 158 3 161 9
rect 212 3 215 9
rect -94 0 251 3
rect 74 -3 79 0
rect 180 -3 184 0
rect 6 -6 255 -3
rect 6 -11 9 -6
rect 52 -12 55 -6
rect 106 -12 109 -6
rect 162 -12 165 -6
rect 216 -12 219 -6
rect 40 -23 43 -15
rect 40 -27 41 -23
rect 23 -36 26 -33
rect 40 -49 43 -27
rect 86 -29 89 -16
rect 86 -32 96 -29
rect 128 -32 131 -28
rect 140 -26 143 -16
rect 140 -29 159 -26
rect 188 -26 191 -25
rect 55 -36 57 -33
rect 77 -36 78 -33
rect 86 -41 89 -32
rect 53 -44 89 -41
rect 53 -49 56 -44
rect 86 -49 89 -44
rect 93 -41 96 -32
rect 107 -36 111 -34
rect 128 -35 132 -32
rect 107 -37 114 -36
rect 140 -41 143 -29
rect 190 -30 191 -26
rect 188 -32 191 -30
rect 164 -36 167 -33
rect 196 -36 199 -16
rect 222 -23 223 -19
rect 220 -32 223 -23
rect 250 -27 253 -16
rect 220 -35 221 -32
rect 239 -36 242 -34
rect 239 -37 245 -36
rect 196 -41 199 -40
rect 250 -41 253 -31
rect 107 -44 143 -41
rect 107 -49 110 -44
rect 140 -49 143 -44
rect 163 -44 199 -41
rect 163 -49 166 -44
rect 196 -49 199 -44
rect 217 -44 253 -41
rect 217 -49 220 -44
rect 250 -49 253 -44
rect 6 -72 9 -53
rect 69 -72 72 -53
rect 79 -72 82 -67
rect 123 -72 126 -53
rect 133 -72 136 -67
rect 179 -72 182 -53
rect 189 -72 192 -67
rect 233 -72 236 -53
rect 243 -72 246 -67
rect 264 -72 269 69
rect 4 -75 269 -72
<< metal2 >>
rect -7 41 73 44
rect -7 35 -4 41
rect -46 32 -4 35
rect 69 34 72 41
rect 93 39 152 42
rect 26 31 47 34
rect 73 31 99 34
rect 103 31 104 34
rect 149 33 152 39
rect 173 34 192 37
rect 149 30 156 33
rect 173 29 176 34
rect 196 35 235 36
rect 196 33 231 35
rect -31 21 -19 24
rect -22 -43 -19 21
rect 41 21 123 24
rect 186 24 245 27
rect 156 19 159 22
rect 156 16 214 19
rect 145 -3 149 15
rect 26 -7 149 -3
rect 26 -33 30 -7
rect 145 -8 149 -7
rect 160 -22 218 -19
rect 45 -27 127 -24
rect 160 -25 163 -22
rect 190 -30 249 -27
rect 30 -37 51 -34
rect 77 -37 103 -34
rect 107 -37 108 -34
rect 153 -36 160 -33
rect 73 -43 76 -37
rect -22 -46 76 -43
rect 153 -42 156 -36
rect 200 -38 235 -36
rect 200 -39 239 -38
rect 97 -45 156 -42
<< ntransistor >>
rect -55 9 -53 12
rect 17 8 19 11
rect 56 8 58 14
rect 77 8 79 14
rect 110 8 112 14
rect 131 8 133 14
rect 166 8 168 14
rect 187 8 189 14
rect 220 8 222 14
rect 241 8 243 14
rect 21 -14 23 -11
rect 60 -17 62 -11
rect 81 -17 83 -11
rect 114 -17 116 -11
rect 135 -17 137 -11
rect 170 -17 172 -11
rect 191 -17 193 -11
rect 224 -17 226 -11
rect 245 -17 247 -11
<< ptransistor >>
rect -55 45 -53 51
rect 17 45 19 51
rect 56 45 58 51
rect 77 45 79 51
rect 110 45 112 51
rect 131 45 133 51
rect 166 45 168 51
rect 187 45 189 51
rect 220 45 222 51
rect 241 45 243 51
rect 21 -54 23 -48
rect 60 -54 62 -48
rect 81 -54 83 -48
rect 114 -54 116 -48
rect 135 -54 137 -48
rect 170 -54 172 -48
rect 191 -54 193 -48
rect 224 -54 226 -48
rect 245 -54 247 -48
<< polycontact >>
rect -57 30 -53 34
rect 15 29 19 33
rect 53 29 57 33
rect 74 29 78 33
rect 107 29 111 33
rect 128 29 132 33
rect 163 29 167 33
rect 184 29 188 33
rect 217 29 221 33
rect 238 29 242 33
rect 19 -36 23 -32
rect 57 -36 61 -32
rect 78 -36 82 -32
rect 111 -36 115 -32
rect 132 -36 136 -32
rect 167 -36 171 -32
rect 188 -36 192 -32
rect 221 -36 225 -32
rect 242 -36 246 -32
<< ndcontact >>
rect -70 9 -66 13
rect -36 9 -32 13
rect 2 8 6 12
rect 36 8 40 12
rect 48 9 52 13
rect 82 9 86 13
rect 102 9 106 13
rect 136 9 140 13
rect 158 9 162 13
rect 192 9 196 13
rect 212 9 216 13
rect 246 9 250 13
rect 6 -15 10 -11
rect 40 -15 44 -11
rect 52 -16 56 -12
rect 86 -16 90 -12
rect 106 -16 110 -12
rect 140 -16 144 -12
rect 162 -16 166 -12
rect 196 -16 200 -12
rect 216 -16 220 -12
rect 250 -16 254 -12
<< pdcontact >>
rect -81 46 -77 50
rect -37 46 -31 52
rect 2 46 6 50
rect 35 46 39 50
rect 48 46 52 50
rect 65 46 69 50
rect 82 46 86 50
rect 102 46 106 50
rect 119 46 123 50
rect 136 46 140 50
rect 158 46 162 50
rect 175 46 179 50
rect 192 46 196 50
rect 212 46 216 50
rect 229 46 233 50
rect 246 46 250 50
rect 6 -53 10 -49
rect 39 -53 43 -49
rect 52 -53 56 -49
rect 69 -53 73 -49
rect 86 -53 90 -49
rect 106 -53 110 -49
rect 123 -53 127 -49
rect 140 -53 144 -49
rect 162 -53 166 -49
rect 179 -53 183 -49
rect 196 -53 200 -49
rect 216 -53 220 -49
rect 233 -53 237 -49
rect 250 -53 254 -49
<< m2contact >>
rect -50 31 -46 35
rect 22 30 26 34
rect -35 21 -31 25
rect 47 30 51 34
rect 69 30 73 34
rect 89 38 93 42
rect 99 30 103 34
rect 37 20 41 24
rect 123 21 127 25
rect 156 30 160 34
rect 192 33 196 37
rect 155 22 159 26
rect 172 25 176 29
rect 182 23 186 27
rect 145 15 149 19
rect 231 31 235 35
rect 245 24 249 28
rect 214 16 218 20
rect 41 -27 45 -23
rect 26 -37 30 -33
rect 127 -28 131 -24
rect 159 -29 163 -25
rect 51 -37 55 -33
rect 73 -37 77 -33
rect 103 -37 107 -33
rect 186 -30 190 -26
rect 160 -37 164 -33
rect 218 -23 222 -19
rect 249 -31 253 -27
rect 196 -40 200 -36
rect 235 -38 239 -34
rect 93 -45 97 -41
<< nsubstratencontact >>
rect 75 60 79 64
rect 129 60 133 64
rect 185 60 189 64
rect 239 60 243 64
rect 79 -67 83 -63
rect 133 -67 137 -63
rect 189 -67 193 -63
rect 243 -67 247 -63
<< labels >>
rlabel metal1 231 1 231 1 1 gnd
rlabel polycontact 55 31 55 31 1 D
rlabel metal1 37 30 37 30 1 D_bar
rlabel polycontact 76 31 76 31 1 en
rlabel ndiffusion 65 11 65 11 1 n1
rlabel ndiffusion 121 11 121 11 1 n2
rlabel ndiffusion 177 11 177 11 1 n3
rlabel ndiffusion 231 11 231 11 1 n4
rlabel metal1 139 24 139 24 1 out_n2
rlabel metal1 84 28 84 28 1 out_n1
rlabel m2contact 198 -38 198 -38 5 q
rlabel m2contact 252 -30 252 -30 7 q_bar
rlabel metal1 235 -73 235 -73 1 vdd
rlabel metal1 235 -4 235 -4 5 gnd
rlabel m2contact -34 23 -34 23 1 en_bar
rlabel polycontact 59 -34 59 -34 1 q_l1
rlabel m2contact 248 27 248 27 1 q_l1_bar
rlabel ndiffusion 235 -14 235 -14 1 n10
rlabel ndiffusion 181 -14 181 -14 1 n9
rlabel ndiffusion 125 -14 125 -14 1 n8
rlabel metal1 143 -27 143 -27 1 out_n8
rlabel metal1 88 -31 88 -31 1 out_n7
rlabel ndiffusion 69 -14 69 -14 1 n7
rlabel metal1 41 -30 41 -30 1 n6
<< end >>
