magic
tech scmos
timestamp 1521568401
<< pwell >>
rect 0 0 104 36
rect 119 0 279 36
<< nwell >>
rect 0 36 104 80
rect 119 36 279 80
<< polysilicon >>
rect 13 70 15 74
rect 36 67 38 72
rect 43 67 45 72
rect 61 70 63 74
rect 71 70 73 74
rect 81 70 83 74
rect 132 70 134 74
rect 26 58 28 63
rect 13 32 15 45
rect 26 42 28 45
rect 155 67 157 72
rect 162 67 164 72
rect 180 70 182 74
rect 190 70 192 74
rect 200 70 202 74
rect 145 58 147 63
rect 19 41 28 42
rect 19 37 20 41
rect 24 40 28 41
rect 24 37 25 40
rect 36 39 38 42
rect 43 39 45 42
rect 61 39 63 42
rect 71 39 73 42
rect 81 39 83 42
rect 19 36 25 37
rect 13 31 19 32
rect 13 27 14 31
rect 18 27 19 31
rect 13 26 19 27
rect 13 23 15 26
rect 23 23 25 36
rect 33 38 39 39
rect 33 34 34 38
rect 38 34 39 38
rect 33 33 39 34
rect 43 38 65 39
rect 43 34 53 38
rect 57 34 60 38
rect 64 34 65 38
rect 43 33 65 34
rect 69 38 75 39
rect 69 34 70 38
rect 74 34 75 38
rect 69 33 75 34
rect 79 38 85 39
rect 79 34 80 38
rect 84 34 85 38
rect 79 33 85 34
rect 33 30 35 33
rect 43 30 45 33
rect 63 30 65 33
rect 70 30 72 33
rect 13 6 15 10
rect 23 8 25 13
rect 33 11 35 16
rect 43 11 45 16
rect 81 24 83 33
rect 132 32 134 45
rect 145 42 147 45
rect 257 70 259 74
rect 264 70 266 74
rect 244 60 246 65
rect 138 41 147 42
rect 138 37 139 41
rect 143 40 147 41
rect 143 37 144 40
rect 155 39 157 42
rect 162 39 164 42
rect 180 39 182 42
rect 190 39 192 42
rect 200 39 202 42
rect 244 39 246 42
rect 257 39 259 49
rect 264 46 266 49
rect 264 45 270 46
rect 264 41 265 45
rect 269 41 270 45
rect 264 40 270 41
rect 138 36 144 37
rect 132 31 138 32
rect 132 27 133 31
rect 137 27 138 31
rect 132 26 138 27
rect 132 23 134 26
rect 142 23 144 36
rect 152 38 158 39
rect 152 34 153 38
rect 157 34 158 38
rect 152 33 158 34
rect 162 38 184 39
rect 162 34 172 38
rect 176 34 179 38
rect 183 34 184 38
rect 162 33 184 34
rect 188 38 194 39
rect 188 34 189 38
rect 193 34 194 38
rect 188 33 194 34
rect 198 38 204 39
rect 198 34 199 38
rect 203 34 204 38
rect 198 33 204 34
rect 244 38 250 39
rect 244 34 245 38
rect 249 34 250 38
rect 244 33 250 34
rect 254 38 260 39
rect 254 34 255 38
rect 259 34 260 38
rect 254 33 260 34
rect 152 30 154 33
rect 162 30 164 33
rect 182 30 184 33
rect 189 30 191 33
rect 63 6 65 10
rect 70 6 72 10
rect 81 6 83 10
rect 132 6 134 10
rect 142 8 144 13
rect 152 11 154 16
rect 162 11 164 16
rect 200 24 202 33
rect 244 30 246 33
rect 254 30 256 33
rect 264 30 266 40
rect 244 16 246 21
rect 254 19 256 24
rect 264 19 266 24
rect 182 6 184 10
rect 189 6 191 10
rect 200 6 202 10
<< ndiffusion >>
rect 28 23 33 30
rect 6 22 13 23
rect 6 18 7 22
rect 11 18 13 22
rect 6 17 13 18
rect 8 10 13 17
rect 15 18 23 23
rect 15 14 17 18
rect 21 14 23 18
rect 15 13 23 14
rect 25 21 33 23
rect 25 17 27 21
rect 31 17 33 21
rect 25 16 33 17
rect 35 29 43 30
rect 35 25 37 29
rect 41 25 43 29
rect 35 16 43 25
rect 45 29 52 30
rect 45 25 47 29
rect 51 25 52 29
rect 45 22 52 25
rect 58 23 63 30
rect 45 18 47 22
rect 51 18 52 22
rect 45 16 52 18
rect 56 22 63 23
rect 56 18 57 22
rect 61 18 63 22
rect 56 17 63 18
rect 25 13 30 16
rect 15 10 20 13
rect 58 10 63 17
rect 65 10 70 30
rect 72 24 79 30
rect 72 15 81 24
rect 72 11 74 15
rect 78 11 81 15
rect 72 10 81 11
rect 83 22 90 24
rect 147 23 152 30
rect 83 18 85 22
rect 89 18 90 22
rect 83 17 90 18
rect 125 22 132 23
rect 125 18 126 22
rect 130 18 132 22
rect 125 17 132 18
rect 83 10 88 17
rect 127 10 132 17
rect 134 18 142 23
rect 134 14 136 18
rect 140 14 142 18
rect 134 13 142 14
rect 144 21 152 23
rect 144 17 146 21
rect 150 17 152 21
rect 144 16 152 17
rect 154 29 162 30
rect 154 25 156 29
rect 160 25 162 29
rect 154 16 162 25
rect 164 29 171 30
rect 164 25 166 29
rect 170 25 171 29
rect 164 22 171 25
rect 177 23 182 30
rect 164 18 166 22
rect 170 18 171 22
rect 164 16 171 18
rect 175 22 182 23
rect 175 18 176 22
rect 180 18 182 22
rect 175 17 182 18
rect 144 13 149 16
rect 134 10 139 13
rect 177 10 182 17
rect 184 10 189 30
rect 191 24 198 30
rect 237 29 244 30
rect 237 25 238 29
rect 242 25 244 29
rect 237 24 244 25
rect 191 15 200 24
rect 191 11 193 15
rect 197 11 200 15
rect 191 10 200 11
rect 202 22 209 24
rect 202 18 204 22
rect 208 18 209 22
rect 239 21 244 24
rect 246 24 254 30
rect 256 29 264 30
rect 256 25 258 29
rect 262 25 264 29
rect 256 24 264 25
rect 266 24 273 30
rect 246 21 252 24
rect 202 17 209 18
rect 202 10 207 17
rect 248 17 252 21
rect 268 17 273 24
rect 248 16 254 17
rect 248 12 249 16
rect 253 12 254 16
rect 248 11 254 12
rect 267 16 273 17
rect 267 12 268 16
rect 272 12 273 16
rect 267 11 273 12
<< pdiffusion >>
rect 8 58 13 70
rect 6 57 13 58
rect 6 53 7 57
rect 11 53 13 57
rect 6 50 13 53
rect 6 46 7 50
rect 11 46 13 50
rect 6 45 13 46
rect 15 69 24 70
rect 15 65 18 69
rect 22 65 24 69
rect 47 69 61 70
rect 47 67 53 69
rect 15 58 24 65
rect 31 58 36 67
rect 15 45 26 58
rect 28 50 36 58
rect 28 46 30 50
rect 34 46 36 50
rect 28 45 36 46
rect 31 42 36 45
rect 38 42 43 67
rect 45 65 53 67
rect 57 65 61 69
rect 45 62 61 65
rect 45 58 53 62
rect 57 58 61 62
rect 45 42 61 58
rect 63 61 71 70
rect 63 57 65 61
rect 69 57 71 61
rect 63 54 71 57
rect 63 50 65 54
rect 69 50 71 54
rect 63 42 71 50
rect 73 69 81 70
rect 73 65 75 69
rect 79 65 81 69
rect 73 62 81 65
rect 73 58 75 62
rect 79 58 81 62
rect 73 42 81 58
rect 83 55 88 70
rect 127 58 132 70
rect 125 57 132 58
rect 83 54 90 55
rect 83 50 85 54
rect 89 50 90 54
rect 83 47 90 50
rect 83 43 85 47
rect 89 43 90 47
rect 125 53 126 57
rect 130 53 132 57
rect 125 50 132 53
rect 125 46 126 50
rect 130 46 132 50
rect 125 45 132 46
rect 134 69 143 70
rect 134 65 137 69
rect 141 65 143 69
rect 166 69 180 70
rect 166 67 172 69
rect 134 58 143 65
rect 150 58 155 67
rect 134 45 145 58
rect 147 50 155 58
rect 147 46 149 50
rect 153 46 155 50
rect 147 45 155 46
rect 83 42 90 43
rect 150 42 155 45
rect 157 42 162 67
rect 164 65 172 67
rect 176 65 180 69
rect 164 62 180 65
rect 164 58 172 62
rect 176 58 180 62
rect 164 42 180 58
rect 182 61 190 70
rect 182 57 184 61
rect 188 57 190 61
rect 182 54 190 57
rect 182 50 184 54
rect 188 50 190 54
rect 182 42 190 50
rect 192 69 200 70
rect 192 65 194 69
rect 198 65 200 69
rect 192 62 200 65
rect 192 58 194 62
rect 198 58 200 62
rect 192 42 200 58
rect 202 55 207 70
rect 248 69 257 70
rect 248 65 249 69
rect 253 65 257 69
rect 248 60 257 65
rect 237 59 244 60
rect 237 55 238 59
rect 242 55 244 59
rect 202 54 209 55
rect 202 50 204 54
rect 208 50 209 54
rect 202 47 209 50
rect 237 52 244 55
rect 237 48 238 52
rect 242 48 244 52
rect 237 47 244 48
rect 202 43 204 47
rect 208 43 209 47
rect 202 42 209 43
rect 239 42 244 47
rect 246 49 257 60
rect 259 49 264 70
rect 266 63 271 70
rect 266 62 273 63
rect 266 58 268 62
rect 272 58 273 62
rect 266 57 273 58
rect 266 49 271 57
rect 246 42 254 49
<< metal1 >>
rect 2 72 277 76
rect 2 69 239 72
rect 2 68 18 69
rect 17 65 18 68
rect 22 68 53 69
rect 22 65 23 68
rect 52 65 53 68
rect 57 68 75 69
rect 57 65 58 68
rect 52 62 58 65
rect 74 65 75 68
rect 79 68 137 69
rect 79 65 80 68
rect 136 65 137 68
rect 141 68 172 69
rect 141 65 142 68
rect 171 65 172 68
rect 176 68 194 69
rect 176 65 177 68
rect 74 62 80 65
rect 171 62 177 65
rect 193 65 194 68
rect 198 68 239 69
rect 243 69 277 72
rect 243 68 249 69
rect 198 65 199 68
rect 248 65 249 68
rect 253 68 277 69
rect 253 65 254 68
rect 193 62 199 65
rect 6 58 19 62
rect 52 58 53 62
rect 57 58 58 62
rect 65 61 69 62
rect 6 57 11 58
rect 6 53 7 57
rect 22 54 46 58
rect 74 58 75 62
rect 79 58 80 62
rect 125 58 138 62
rect 171 58 172 62
rect 176 58 177 62
rect 184 61 188 62
rect 65 54 69 57
rect 125 57 130 58
rect 85 54 91 55
rect 6 50 11 53
rect 6 46 7 50
rect 6 45 11 46
rect 20 50 26 54
rect 30 50 34 51
rect 42 50 65 54
rect 69 50 82 54
rect 6 37 10 45
rect 20 41 24 50
rect 20 36 24 37
rect 27 42 34 46
rect 37 42 75 46
rect 6 23 10 33
rect 27 31 31 42
rect 37 39 42 42
rect 34 38 42 39
rect 70 38 74 42
rect 38 34 42 38
rect 52 34 53 38
rect 57 34 60 38
rect 64 34 67 38
rect 34 33 42 34
rect 13 27 14 31
rect 18 29 31 31
rect 47 29 51 30
rect 18 27 37 29
rect 27 25 37 27
rect 41 25 42 29
rect 54 25 58 34
rect 70 33 74 34
rect 78 39 82 50
rect 89 52 91 54
rect 125 53 126 57
rect 141 54 165 58
rect 193 58 194 62
rect 198 58 199 62
rect 237 62 241 63
rect 237 59 250 62
rect 184 54 188 57
rect 237 55 238 59
rect 242 58 250 59
rect 256 58 268 62
rect 272 58 273 62
rect 204 54 210 55
rect 89 50 105 52
rect 85 49 105 50
rect 125 50 130 53
rect 85 47 91 49
rect 89 43 91 47
rect 85 42 91 43
rect 78 38 84 39
rect 78 34 80 38
rect 78 33 84 34
rect 78 30 82 33
rect 62 26 82 30
rect 6 22 11 23
rect 6 18 7 22
rect 47 22 51 25
rect 62 22 66 26
rect 87 22 91 42
rect 6 17 11 18
rect 17 18 21 19
rect 26 17 27 21
rect 31 18 47 21
rect 56 18 57 22
rect 61 18 66 22
rect 69 18 85 22
rect 89 18 91 22
rect 125 46 126 50
rect 125 45 130 46
rect 139 50 145 54
rect 149 50 153 51
rect 161 50 184 54
rect 188 50 201 54
rect 125 23 129 45
rect 139 41 143 50
rect 139 36 143 37
rect 146 42 153 46
rect 156 42 194 46
rect 146 31 150 42
rect 156 39 161 42
rect 153 38 161 39
rect 189 38 193 42
rect 157 34 161 38
rect 169 34 172 38
rect 176 34 179 38
rect 183 34 186 38
rect 153 33 161 34
rect 132 27 133 31
rect 137 29 150 31
rect 166 29 170 30
rect 137 27 156 29
rect 146 25 156 27
rect 160 25 161 29
rect 173 25 177 34
rect 189 33 193 34
rect 197 39 201 50
rect 208 50 210 54
rect 204 47 210 50
rect 208 43 210 47
rect 204 42 210 43
rect 197 38 203 39
rect 197 34 199 38
rect 197 33 203 34
rect 206 38 210 42
rect 197 30 201 33
rect 181 26 201 30
rect 125 22 130 23
rect 125 18 126 22
rect 166 22 170 25
rect 181 22 185 26
rect 206 22 210 34
rect 237 52 242 55
rect 256 54 260 58
rect 237 48 238 52
rect 237 47 242 48
rect 245 50 260 54
rect 269 53 273 55
rect 237 30 241 47
rect 245 38 249 50
rect 269 49 272 53
rect 269 46 273 49
rect 252 45 273 46
rect 252 42 265 45
rect 264 41 265 42
rect 269 42 273 45
rect 269 41 270 42
rect 252 34 255 38
rect 259 34 272 38
rect 237 29 242 30
rect 237 25 238 29
rect 245 29 249 34
rect 245 25 258 29
rect 262 25 263 29
rect 269 25 273 34
rect 237 24 242 25
rect 31 17 51 18
rect 125 17 130 18
rect 136 18 140 19
rect 17 12 21 14
rect 73 12 74 15
rect 2 11 74 12
rect 78 12 79 15
rect 145 17 146 21
rect 150 18 166 21
rect 175 18 176 22
rect 180 18 185 22
rect 188 18 204 22
rect 208 18 210 22
rect 150 17 170 18
rect 136 12 140 14
rect 192 12 193 15
rect 78 11 193 12
rect 197 12 198 15
rect 248 12 249 16
rect 253 12 254 16
rect 267 12 268 16
rect 272 12 273 16
rect 197 11 239 12
rect 2 8 239 11
rect 243 8 277 12
rect 2 4 277 8
<< metal2 >>
rect 109 49 272 52
rect -1 34 6 37
rect 10 34 165 37
rect 210 34 272 37
<< ntransistor >>
rect 13 10 15 23
rect 23 13 25 23
rect 33 16 35 30
rect 43 16 45 30
rect 63 10 65 30
rect 70 10 72 30
rect 81 10 83 24
rect 132 10 134 23
rect 142 13 144 23
rect 152 16 154 30
rect 162 16 164 30
rect 182 10 184 30
rect 189 10 191 30
rect 200 10 202 24
rect 244 21 246 30
rect 254 24 256 30
rect 264 24 266 30
<< ptransistor >>
rect 13 45 15 70
rect 26 45 28 58
rect 36 42 38 67
rect 43 42 45 67
rect 61 42 63 70
rect 71 42 73 70
rect 81 42 83 70
rect 132 45 134 70
rect 145 45 147 58
rect 155 42 157 67
rect 162 42 164 67
rect 180 42 182 70
rect 190 42 192 70
rect 200 42 202 70
rect 244 42 246 60
rect 257 49 259 70
rect 264 49 266 70
<< polycontact >>
rect 20 37 24 41
rect 14 27 18 31
rect 34 34 38 38
rect 53 34 57 38
rect 60 34 64 38
rect 70 34 74 38
rect 80 34 84 38
rect 139 37 143 41
rect 265 41 269 45
rect 133 27 137 31
rect 153 34 157 38
rect 172 34 176 38
rect 179 34 183 38
rect 189 34 193 38
rect 199 34 203 38
rect 245 34 249 38
rect 255 34 259 38
<< ndcontact >>
rect 7 18 11 22
rect 17 14 21 18
rect 27 17 31 21
rect 37 25 41 29
rect 47 25 51 29
rect 47 18 51 22
rect 57 18 61 22
rect 74 11 78 15
rect 85 18 89 22
rect 126 18 130 22
rect 136 14 140 18
rect 146 17 150 21
rect 156 25 160 29
rect 166 25 170 29
rect 166 18 170 22
rect 176 18 180 22
rect 238 25 242 29
rect 193 11 197 15
rect 204 18 208 22
rect 258 25 262 29
rect 249 12 253 16
rect 268 12 272 16
<< pdcontact >>
rect 7 53 11 57
rect 7 46 11 50
rect 18 65 22 69
rect 30 46 34 50
rect 53 65 57 69
rect 53 58 57 62
rect 65 57 69 61
rect 65 50 69 54
rect 75 65 79 69
rect 75 58 79 62
rect 85 50 89 54
rect 85 43 89 47
rect 126 53 130 57
rect 126 46 130 50
rect 137 65 141 69
rect 149 46 153 50
rect 172 65 176 69
rect 172 58 176 62
rect 184 57 188 61
rect 184 50 188 54
rect 194 65 198 69
rect 194 58 198 62
rect 249 65 253 69
rect 238 55 242 59
rect 204 50 208 54
rect 238 48 242 52
rect 204 43 208 47
rect 268 58 272 62
<< m2contact >>
rect 6 33 10 37
rect 105 49 109 53
rect 165 34 169 38
rect 206 34 210 38
rect 272 49 276 53
rect 272 34 276 38
<< psubstratepcontact >>
rect 239 8 243 12
<< nsubstratencontact >>
rect 239 68 243 72
<< psubstratepdiff >>
rect 238 12 244 13
rect 238 8 239 12
rect 243 8 244 12
rect 238 7 244 8
<< nsubstratendiff >>
rect 238 72 244 73
rect 238 68 239 72
rect 243 68 244 72
rect 238 67 244 68
<< labels >>
rlabel polycontact 16 29 16 29 6 son
rlabel polycontact 22 39 22 39 6 con
rlabel polysilicon 82 40 82 40 6 con
rlabel metal1 16 60 16 60 6 so
rlabel metal1 22 29 22 29 6 son
rlabel metal1 32 46 32 46 6 son
rlabel metal1 22 45 22 45 6 con
rlabel metal1 52 8 52 8 6 vss
rlabel metal1 49 23 49 23 6 n2
rlabel metal1 38 19 38 19 6 n2
rlabel metal1 34 27 34 27 6 son
rlabel metal1 56 32 56 32 6 a
rlabel metal1 40 40 40 40 6 b
rlabel metal1 56 44 56 44 6 b
rlabel metal1 48 44 48 44 6 b
rlabel metal1 52 72 52 72 6 vdd
rlabel metal1 72 20 72 20 6 co
rlabel metal1 80 20 80 20 6 co
rlabel metal1 61 20 61 20 6 con
rlabel metal1 64 36 64 36 6 a
rlabel metal1 64 44 64 44 6 b
rlabel metal1 72 44 72 44 6 b
rlabel metal1 80 40 80 40 6 con
rlabel metal1 62 52 62 52 6 con
rlabel metal1 67 56 67 56 6 con
rlabel ndcontact 88 20 88 20 6 co
rlabel metal1 88 48 88 48 6 co
rlabel polycontact 135 29 135 29 6 son
rlabel polycontact 141 39 141 39 6 con
rlabel polysilicon 201 40 201 40 6 con
rlabel metal1 141 29 141 29 6 son
rlabel metal1 151 46 151 46 6 son
rlabel metal1 141 45 141 45 6 con
rlabel metal1 171 8 171 8 6 vss
rlabel metal1 168 23 168 23 6 n2
rlabel metal1 157 19 157 19 6 n2
rlabel metal1 153 27 153 27 6 son
rlabel metal1 171 72 171 72 6 vdd
rlabel metal1 180 20 180 20 6 con
rlabel metal1 199 40 199 40 6 con
rlabel metal1 181 52 181 52 6 con
rlabel metal1 186 56 186 56 6 con
rlabel metal1 175 44 175 44 1 c
rlabel metal1 207 48 207 48 1 c1
rlabel polycontact 247 36 247 36 6 zn
rlabel metal1 247 39 247 39 6 zn
rlabel metal1 255 8 255 8 6 vss
rlabel metal1 254 27 254 27 6 zn
rlabel metal1 255 72 255 72 6 vdd
rlabel metal1 264 60 264 60 6 zn
rlabel metal1 238 42 238 42 1 carry
rlabel metal1 127 40 127 40 1 sum
rlabel metal1 8 42 8 42 1 so
<< end >>
