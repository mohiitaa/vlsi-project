magic
tech scmos
timestamp 1522987514
<< nwell >>
rect 6 113 185 139
rect 198 113 239 139
rect 254 113 295 139
rect 308 113 349 139
rect 102 8 189 34
rect 202 8 243 34
rect 258 8 299 34
rect 312 8 353 34
<< polysilicon >>
rect 43 126 45 128
rect 115 126 117 132
rect 154 126 156 132
rect 175 126 177 132
rect 208 126 210 132
rect 229 126 231 132
rect 264 126 266 132
rect 285 126 287 132
rect 318 126 320 132
rect 339 126 341 132
rect 43 109 45 120
rect 115 108 117 120
rect 154 108 156 120
rect 175 108 177 120
rect 208 108 210 120
rect 229 108 231 120
rect 264 108 266 120
rect 285 108 287 120
rect 318 108 320 120
rect 339 108 341 120
rect 43 87 45 105
rect 155 104 156 108
rect 176 104 177 108
rect 209 104 210 108
rect 230 104 231 108
rect 265 104 266 108
rect 286 104 287 108
rect 319 104 320 108
rect 340 104 341 108
rect 43 81 45 84
rect 115 86 117 104
rect 154 89 156 104
rect 175 89 177 104
rect 208 89 210 104
rect 229 89 231 104
rect 264 89 266 104
rect 285 89 287 104
rect 318 89 320 104
rect 339 89 341 104
rect 115 80 117 83
rect 154 80 156 83
rect 175 80 177 83
rect 208 80 210 83
rect 229 80 231 83
rect 264 80 266 83
rect 285 80 287 83
rect 318 80 320 83
rect 339 80 341 83
rect 119 64 121 67
rect 158 64 160 67
rect 179 64 181 67
rect 212 64 214 67
rect 233 64 235 67
rect 268 64 270 67
rect 289 64 291 67
rect 322 64 324 67
rect 343 64 345 67
rect 119 43 121 61
rect 158 43 160 58
rect 179 43 181 58
rect 212 43 214 58
rect 233 43 235 58
rect 268 43 270 58
rect 289 43 291 58
rect 322 43 324 58
rect 343 43 345 58
rect 159 39 160 43
rect 180 39 181 43
rect 213 39 214 43
rect 234 39 235 43
rect 269 39 270 43
rect 290 39 291 43
rect 323 39 324 43
rect 344 39 345 43
rect 119 27 121 39
rect 158 27 160 39
rect 179 27 181 39
rect 212 27 214 39
rect 233 27 235 39
rect 268 27 270 39
rect 289 27 291 39
rect 322 27 324 39
rect 343 27 345 39
rect 119 15 121 21
rect 158 15 160 21
rect 179 15 181 21
rect 212 15 214 21
rect 233 15 235 21
rect 268 15 270 21
rect 289 15 291 21
rect 322 15 324 21
rect 343 15 345 21
<< ndiffusion >>
rect 32 84 43 87
rect 45 84 62 87
rect 144 88 154 89
rect 104 83 115 86
rect 117 83 134 86
rect 144 84 146 88
rect 150 84 154 88
rect 144 83 154 84
rect 156 83 175 89
rect 177 88 185 89
rect 177 84 180 88
rect 184 84 185 88
rect 177 83 185 84
rect 198 88 208 89
rect 198 84 200 88
rect 204 84 208 88
rect 198 83 208 84
rect 210 83 229 89
rect 231 88 239 89
rect 231 84 234 88
rect 238 84 239 88
rect 231 83 239 84
rect 254 88 264 89
rect 254 84 256 88
rect 260 84 264 88
rect 254 83 264 84
rect 266 83 285 89
rect 287 88 295 89
rect 287 84 290 88
rect 294 84 295 88
rect 287 83 295 84
rect 308 88 318 89
rect 308 84 310 88
rect 314 84 318 88
rect 308 83 318 84
rect 320 83 339 89
rect 341 88 349 89
rect 341 84 344 88
rect 348 84 349 88
rect 341 83 349 84
rect 108 61 119 64
rect 121 61 138 64
rect 148 63 158 64
rect 148 59 150 63
rect 154 59 158 63
rect 148 58 158 59
rect 160 58 179 64
rect 181 63 189 64
rect 181 59 184 63
rect 188 59 189 63
rect 181 58 189 59
rect 202 63 212 64
rect 202 59 204 63
rect 208 59 212 63
rect 202 58 212 59
rect 214 58 233 64
rect 235 63 243 64
rect 235 59 238 63
rect 242 59 243 63
rect 235 58 243 59
rect 258 63 268 64
rect 258 59 260 63
rect 264 59 268 63
rect 258 58 268 59
rect 270 58 289 64
rect 291 63 299 64
rect 291 59 294 63
rect 298 59 299 63
rect 291 58 299 59
rect 312 63 322 64
rect 312 59 314 63
rect 318 59 322 63
rect 312 58 322 59
rect 324 58 343 64
rect 345 63 353 64
rect 345 59 348 63
rect 352 59 353 63
rect 345 58 353 59
<< pdiffusion >>
rect 12 125 43 126
rect 12 121 17 125
rect 21 121 43 125
rect 12 120 43 121
rect 45 121 61 126
rect 67 121 80 126
rect 45 120 80 121
rect 100 125 115 126
rect 104 121 115 125
rect 100 120 115 121
rect 117 125 137 126
rect 117 121 133 125
rect 117 120 137 121
rect 144 125 154 126
rect 144 121 146 125
rect 150 121 154 125
rect 144 120 154 121
rect 156 125 175 126
rect 156 121 163 125
rect 167 121 175 125
rect 156 120 175 121
rect 177 125 185 126
rect 177 121 180 125
rect 184 121 185 125
rect 177 120 185 121
rect 198 125 208 126
rect 198 121 200 125
rect 204 121 208 125
rect 198 120 208 121
rect 210 125 229 126
rect 210 121 217 125
rect 221 121 229 125
rect 210 120 229 121
rect 231 125 239 126
rect 231 121 234 125
rect 238 121 239 125
rect 231 120 239 121
rect 254 125 264 126
rect 254 121 256 125
rect 260 121 264 125
rect 254 120 264 121
rect 266 125 285 126
rect 266 121 273 125
rect 277 121 285 125
rect 266 120 285 121
rect 287 125 295 126
rect 287 121 290 125
rect 294 121 295 125
rect 287 120 295 121
rect 308 125 318 126
rect 308 121 310 125
rect 314 121 318 125
rect 308 120 318 121
rect 320 125 339 126
rect 320 121 327 125
rect 331 121 339 125
rect 320 120 339 121
rect 341 125 349 126
rect 341 121 344 125
rect 348 121 349 125
rect 341 120 349 121
rect 104 26 119 27
rect 108 22 119 26
rect 104 21 119 22
rect 121 26 141 27
rect 121 22 137 26
rect 121 21 141 22
rect 148 26 158 27
rect 148 22 150 26
rect 154 22 158 26
rect 148 21 158 22
rect 160 26 179 27
rect 160 22 167 26
rect 171 22 179 26
rect 160 21 179 22
rect 181 26 189 27
rect 181 22 184 26
rect 188 22 189 26
rect 181 21 189 22
rect 202 26 212 27
rect 202 22 204 26
rect 208 22 212 26
rect 202 21 212 22
rect 214 26 233 27
rect 214 22 221 26
rect 225 22 233 26
rect 214 21 233 22
rect 235 26 243 27
rect 235 22 238 26
rect 242 22 243 26
rect 235 21 243 22
rect 258 26 268 27
rect 258 22 260 26
rect 264 22 268 26
rect 258 21 268 22
rect 270 26 289 27
rect 270 22 277 26
rect 281 22 289 26
rect 270 21 289 22
rect 291 26 299 27
rect 291 22 294 26
rect 298 22 299 26
rect 291 21 299 22
rect 312 26 322 27
rect 312 22 314 26
rect 318 22 322 26
rect 312 21 322 22
rect 324 26 343 27
rect 324 22 331 26
rect 335 22 343 26
rect 324 21 343 22
rect 345 26 353 27
rect 345 22 348 26
rect 352 22 353 26
rect 345 21 353 22
<< metal1 >>
rect 1 144 367 147
rect 17 125 20 144
rect 30 133 84 136
rect 62 127 66 129
rect 62 110 66 121
rect 81 118 84 133
rect 100 125 103 144
rect 163 125 166 144
rect 173 139 176 144
rect 217 125 220 144
rect 227 139 230 144
rect 273 125 276 144
rect 283 139 286 144
rect 327 125 330 144
rect 337 139 340 144
rect 81 115 131 118
rect 45 106 48 109
rect 62 100 65 110
rect 117 105 120 108
rect 62 96 63 100
rect 62 88 65 96
rect 127 95 131 115
rect 134 99 137 121
rect 147 116 150 121
rect 180 116 183 121
rect 147 113 183 116
rect 149 105 151 108
rect 171 105 172 108
rect 180 104 183 113
rect 201 116 204 121
rect 234 116 237 121
rect 201 113 237 116
rect 257 116 260 121
rect 290 116 293 121
rect 257 113 293 116
rect 311 116 314 121
rect 344 116 347 121
rect 311 113 347 116
rect 187 104 190 113
rect 201 108 208 109
rect 201 106 205 108
rect 222 104 226 107
rect 180 101 190 104
rect 134 95 135 99
rect 134 87 137 95
rect 180 88 183 101
rect 222 100 225 104
rect 234 101 237 113
rect 290 112 293 113
rect 258 105 261 108
rect 234 98 253 101
rect 234 88 237 98
rect 282 102 285 104
rect 270 94 273 100
rect 284 98 285 102
rect 282 97 285 98
rect 247 91 273 94
rect 290 88 293 108
rect 314 104 315 107
rect 333 108 339 109
rect 333 106 336 108
rect 314 95 317 104
rect 344 103 347 113
rect 316 91 317 95
rect 344 88 347 99
rect 28 78 31 84
rect 100 78 103 83
rect 146 78 149 84
rect 200 78 203 84
rect 256 78 259 84
rect 310 78 313 84
rect 4 75 349 78
rect 172 72 177 75
rect 278 72 282 75
rect 104 69 353 72
rect 104 64 107 69
rect 150 63 153 69
rect 204 63 207 69
rect 260 63 263 69
rect 314 63 317 69
rect 138 52 141 60
rect 138 48 139 52
rect 121 39 124 42
rect 138 26 141 48
rect 184 46 187 59
rect 184 43 194 46
rect 226 43 229 47
rect 238 49 241 59
rect 238 46 257 49
rect 286 49 289 50
rect 153 39 155 42
rect 175 39 176 42
rect 184 34 187 43
rect 151 31 187 34
rect 151 26 154 31
rect 184 26 187 31
rect 191 34 194 43
rect 205 39 209 41
rect 226 40 230 43
rect 205 38 212 39
rect 238 34 241 46
rect 288 45 289 49
rect 286 43 289 45
rect 262 39 265 42
rect 294 39 297 59
rect 320 52 321 56
rect 318 43 321 52
rect 348 48 351 59
rect 318 40 319 43
rect 337 39 340 41
rect 337 38 343 39
rect 294 34 297 35
rect 348 34 351 44
rect 205 31 241 34
rect 205 26 208 31
rect 238 26 241 31
rect 261 31 297 34
rect 261 26 264 31
rect 294 26 297 31
rect 315 31 351 34
rect 315 26 318 31
rect 348 26 351 31
rect 104 3 107 22
rect 167 3 170 22
rect 177 3 180 8
rect 221 3 224 22
rect 231 3 234 8
rect 277 3 280 22
rect 287 3 290 8
rect 331 3 334 22
rect 341 3 344 8
rect 362 3 367 144
rect 102 0 367 3
<< metal2 >>
rect 1 133 26 136
rect 91 116 171 119
rect 91 110 94 116
rect 52 107 94 110
rect 167 109 170 116
rect 191 114 250 117
rect 124 106 145 109
rect 128 100 131 106
rect 171 106 197 109
rect 201 106 202 109
rect 247 108 250 114
rect 271 109 290 112
rect 247 105 254 108
rect 271 104 274 109
rect 294 110 333 111
rect 294 108 329 110
rect 121 99 131 100
rect 67 96 79 99
rect 121 97 123 99
rect 76 32 79 96
rect 127 97 131 99
rect 139 96 221 99
rect 284 99 343 102
rect 254 94 257 97
rect 254 91 312 94
rect 243 72 247 90
rect 124 68 247 72
rect 124 42 128 68
rect 243 67 247 68
rect 258 53 316 56
rect 143 48 225 51
rect 258 50 261 53
rect 288 45 347 48
rect 128 38 149 41
rect 175 38 201 41
rect 205 38 206 41
rect 251 39 258 42
rect 171 32 174 38
rect 76 29 174 32
rect 251 33 254 39
rect 298 37 333 39
rect 298 36 337 37
rect 195 30 254 33
rect 304 0 307 36
rect 304 -3 402 0
<< ntransistor >>
rect 43 84 45 87
rect 115 83 117 86
rect 154 83 156 89
rect 175 83 177 89
rect 208 83 210 89
rect 229 83 231 89
rect 264 83 266 89
rect 285 83 287 89
rect 318 83 320 89
rect 339 83 341 89
rect 119 61 121 64
rect 158 58 160 64
rect 179 58 181 64
rect 212 58 214 64
rect 233 58 235 64
rect 268 58 270 64
rect 289 58 291 64
rect 322 58 324 64
rect 343 58 345 64
<< ptransistor >>
rect 43 120 45 126
rect 115 120 117 126
rect 154 120 156 126
rect 175 120 177 126
rect 208 120 210 126
rect 229 120 231 126
rect 264 120 266 126
rect 285 120 287 126
rect 318 120 320 126
rect 339 120 341 126
rect 119 21 121 27
rect 158 21 160 27
rect 179 21 181 27
rect 212 21 214 27
rect 233 21 235 27
rect 268 21 270 27
rect 289 21 291 27
rect 322 21 324 27
rect 343 21 345 27
<< polycontact >>
rect 41 105 45 109
rect 113 104 117 108
rect 151 104 155 108
rect 172 104 176 108
rect 205 104 209 108
rect 226 104 230 108
rect 261 104 265 108
rect 282 104 286 108
rect 315 104 319 108
rect 336 104 340 108
rect 117 39 121 43
rect 155 39 159 43
rect 176 39 180 43
rect 209 39 213 43
rect 230 39 234 43
rect 265 39 269 43
rect 286 39 290 43
rect 319 39 323 43
rect 340 39 344 43
<< ndcontact >>
rect 28 84 32 88
rect 62 84 66 88
rect 100 83 104 87
rect 134 83 138 87
rect 146 84 150 88
rect 180 84 184 88
rect 200 84 204 88
rect 234 84 238 88
rect 256 84 260 88
rect 290 84 294 88
rect 310 84 314 88
rect 344 84 348 88
rect 104 60 108 64
rect 138 60 142 64
rect 150 59 154 63
rect 184 59 188 63
rect 204 59 208 63
rect 238 59 242 63
rect 260 59 264 63
rect 294 59 298 63
rect 314 59 318 63
rect 348 59 352 63
<< pdcontact >>
rect 17 121 21 125
rect 61 121 67 127
rect 100 121 104 125
rect 133 121 137 125
rect 146 121 150 125
rect 163 121 167 125
rect 180 121 184 125
rect 200 121 204 125
rect 217 121 221 125
rect 234 121 238 125
rect 256 121 260 125
rect 273 121 277 125
rect 290 121 294 125
rect 310 121 314 125
rect 327 121 331 125
rect 344 121 348 125
rect 104 22 108 26
rect 137 22 141 26
rect 150 22 154 26
rect 167 22 171 26
rect 184 22 188 26
rect 204 22 208 26
rect 221 22 225 26
rect 238 22 242 26
rect 260 22 264 26
rect 277 22 281 26
rect 294 22 298 26
rect 314 22 318 26
rect 331 22 335 26
rect 348 22 352 26
<< m2contact >>
rect 26 133 30 137
rect 48 106 52 110
rect 120 105 124 109
rect 63 96 67 100
rect 123 95 127 99
rect 145 105 149 109
rect 167 105 171 109
rect 187 113 191 117
rect 197 105 201 109
rect 135 95 139 99
rect 221 96 225 100
rect 254 105 258 109
rect 290 108 294 112
rect 253 97 257 101
rect 270 100 274 104
rect 280 98 284 102
rect 243 90 247 94
rect 329 106 333 110
rect 343 99 347 103
rect 312 91 316 95
rect 139 48 143 52
rect 124 38 128 42
rect 225 47 229 51
rect 257 46 261 50
rect 149 38 153 42
rect 171 38 175 42
rect 201 38 205 42
rect 284 45 288 49
rect 258 38 262 42
rect 316 52 320 56
rect 347 44 351 48
rect 294 35 298 39
rect 333 37 337 41
rect 191 30 195 34
<< nsubstratencontact >>
rect 173 135 177 139
rect 227 135 231 139
rect 283 135 287 139
rect 337 135 341 139
rect 177 8 181 12
rect 231 8 235 12
rect 287 8 291 12
rect 341 8 345 12
<< labels >>
rlabel metal1 329 76 329 76 1 gnd
rlabel metal1 333 2 333 2 1 vdd
rlabel metal1 333 71 333 71 5 gnd
rlabel m2contact 64 98 64 98 1 en_bar_D1
rlabel metal1 135 105 135 105 1 D_bar_D1
rlabel polycontact 153 106 153 106 1 D_D1
rlabel polycontact 174 106 174 106 1 en_D1
rlabel metal1 182 103 182 103 1 out_n1_D1
rlabel ndiffusion 163 86 163 86 1 n1_D1
rlabel ndiffusion 219 86 219 86 1 n2_D1
rlabel metal1 237 99 237 99 1 out_n2_D1
rlabel ndiffusion 275 86 275 86 1 n3_D1
rlabel ndiffusion 329 86 329 86 1 n4_D1
rlabel m2contact 346 102 346 102 1 q_l1_bar_D1
rlabel m2contact 350 45 350 45 1 q_bar_D1
rlabel ndiffusion 333 61 333 61 1 n10_D1
rlabel metal1 241 48 241 48 1 out_n8_D1
rlabel ndiffusion 223 61 223 61 1 n8_D1
rlabel metal1 186 44 186 44 1 out_n7_D1
rlabel ndiffusion 167 61 167 61 1 n7_D1
rlabel polycontact 157 41 157 41 1 q_l1_D1
rlabel metal1 139 45 139 45 1 n6_D1
rlabel ndiffusion 279 61 279 61 1 n9_D1
rlabel m2contact 296 37 296 37 1 q_D1
rlabel metal2 399 -2 399 -2 8 q_D1
rlabel metal2 2 135 2 135 3 D_D1
<< end >>
