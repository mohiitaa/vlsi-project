magic
tech scmos
timestamp 1522676175
<< pwell >>
rect 108 233 126 237
rect 106 229 126 233
rect 106 193 154 229
rect 193 193 241 229
rect 286 193 334 229
rect 526 195 574 231
rect 619 195 667 231
rect 706 195 754 231
rect 35 70 178 106
rect 190 70 308 106
rect 364 72 507 108
rect 519 72 637 108
rect 691 75 834 111
rect 846 75 964 111
rect 121 44 169 70
rect 450 46 498 72
rect 777 49 825 75
rect 34 -76 177 -40
rect 189 -76 307 -40
rect 363 -74 506 -38
rect 518 -74 636 -38
rect 690 -71 833 -35
rect 845 -71 963 -35
rect 120 -102 168 -76
rect 449 -100 497 -74
rect 776 -97 824 -71
rect 321 -224 369 -188
rect 414 -224 462 -188
rect 501 -224 549 -188
<< nwell >>
rect 106 150 154 193
rect 193 150 241 193
rect 286 150 334 193
rect 526 158 574 195
rect 619 158 667 195
rect 526 155 667 158
rect 522 152 667 155
rect 706 164 754 195
rect 706 155 767 164
rect 706 152 834 155
rect 35 106 178 150
rect 190 149 334 150
rect 190 106 308 149
rect 364 108 507 152
rect 519 138 834 152
rect 519 108 637 138
rect 691 111 834 138
rect 846 111 964 155
rect 121 37 169 44
rect 450 39 498 46
rect 777 42 825 49
rect 117 24 169 37
rect 446 26 498 39
rect 773 29 825 42
rect 121 8 169 24
rect 450 10 498 26
rect 777 16 825 29
rect 110 4 176 8
rect 440 6 506 10
rect 748 9 859 16
rect 34 -40 177 4
rect 189 -40 307 4
rect 363 -38 506 6
rect 518 -38 636 6
rect 690 0 963 9
rect 690 -35 833 0
rect 845 -35 963 0
rect 120 -109 168 -102
rect 449 -107 497 -100
rect 776 -104 824 -97
rect 116 -122 168 -109
rect 445 -120 497 -107
rect 772 -117 824 -104
rect 120 -146 168 -122
rect 449 -130 497 -120
rect 323 -144 555 -130
rect 776 -141 824 -117
rect 321 -147 555 -144
rect 321 -188 369 -147
rect 414 -188 462 -147
rect 501 -188 549 -147
<< polysilicon >>
rect 119 212 121 217
rect 126 212 128 217
rect 139 210 141 214
rect 206 212 208 217
rect 213 212 215 217
rect 226 210 228 214
rect 299 212 301 217
rect 306 212 308 217
rect 319 210 321 214
rect 539 212 541 216
rect 552 214 554 219
rect 559 214 561 219
rect 632 212 634 216
rect 645 214 647 219
rect 652 214 654 219
rect 719 212 721 216
rect 732 214 734 219
rect 739 214 741 219
rect 119 188 121 201
rect 126 196 128 201
rect 139 196 141 201
rect 125 195 131 196
rect 125 191 126 195
rect 130 191 131 195
rect 125 190 131 191
rect 135 195 141 196
rect 135 191 136 195
rect 140 191 141 195
rect 135 190 141 191
rect 115 187 121 188
rect 115 183 116 187
rect 120 183 121 187
rect 115 182 121 183
rect 119 179 121 182
rect 129 179 131 190
rect 139 186 141 190
rect 206 188 208 201
rect 213 196 215 201
rect 226 196 228 201
rect 212 195 218 196
rect 212 191 213 195
rect 217 191 218 195
rect 212 190 218 191
rect 222 195 228 196
rect 222 191 223 195
rect 227 191 228 195
rect 222 190 228 191
rect 202 187 208 188
rect 202 183 203 187
rect 207 183 208 187
rect 202 182 208 183
rect 206 179 208 182
rect 216 179 218 190
rect 226 186 228 190
rect 299 188 301 201
rect 306 196 308 201
rect 319 196 321 201
rect 305 195 311 196
rect 305 191 306 195
rect 310 191 311 195
rect 305 190 311 191
rect 315 195 321 196
rect 315 191 316 195
rect 320 191 321 195
rect 315 190 321 191
rect 295 187 301 188
rect 119 161 121 166
rect 129 161 131 166
rect 139 164 141 168
rect 295 183 296 187
rect 300 183 301 187
rect 295 182 301 183
rect 299 179 301 182
rect 309 179 311 190
rect 319 186 321 190
rect 539 198 541 203
rect 552 198 554 203
rect 539 197 545 198
rect 539 193 540 197
rect 544 193 545 197
rect 539 192 545 193
rect 549 197 555 198
rect 549 193 550 197
rect 554 193 555 197
rect 549 192 555 193
rect 539 188 541 192
rect 206 161 208 166
rect 216 161 218 166
rect 226 164 228 168
rect 549 181 551 192
rect 559 190 561 203
rect 632 198 634 203
rect 645 198 647 203
rect 632 197 638 198
rect 632 193 633 197
rect 637 193 638 197
rect 632 192 638 193
rect 642 197 648 198
rect 642 193 643 197
rect 647 193 648 197
rect 642 192 648 193
rect 559 189 565 190
rect 559 185 560 189
rect 564 185 565 189
rect 632 188 634 192
rect 559 184 565 185
rect 559 181 561 184
rect 299 161 301 166
rect 309 161 311 166
rect 319 164 321 168
rect 539 166 541 170
rect 642 181 644 192
rect 652 190 654 203
rect 719 198 721 203
rect 732 198 734 203
rect 719 197 725 198
rect 719 193 720 197
rect 724 193 725 197
rect 719 192 725 193
rect 729 197 735 198
rect 729 193 730 197
rect 734 193 735 197
rect 729 192 735 193
rect 652 189 658 190
rect 652 185 653 189
rect 657 185 658 189
rect 719 188 721 192
rect 652 184 658 185
rect 652 181 654 184
rect 549 163 551 168
rect 559 163 561 168
rect 632 166 634 170
rect 729 181 731 192
rect 739 190 741 203
rect 739 189 745 190
rect 739 185 740 189
rect 744 185 745 189
rect 739 184 745 185
rect 739 181 741 184
rect 642 163 644 168
rect 652 163 654 168
rect 719 166 721 170
rect 729 163 731 168
rect 739 163 741 168
rect 127 140 129 144
rect 51 132 57 133
rect 41 124 43 129
rect 51 128 52 132
rect 56 128 57 132
rect 51 127 57 128
rect 51 122 53 127
rect 61 122 63 127
rect 112 124 118 125
rect 112 120 113 124
rect 117 120 118 124
rect 112 119 118 120
rect 41 109 43 112
rect 51 109 53 112
rect 41 108 47 109
rect 41 104 42 108
rect 46 104 47 108
rect 51 106 55 109
rect 41 103 47 104
rect 41 95 43 103
rect 53 92 55 106
rect 61 101 63 112
rect 116 110 118 119
rect 163 140 165 144
rect 211 140 213 144
rect 143 131 145 135
rect 153 131 155 135
rect 196 124 202 125
rect 196 120 197 124
rect 201 120 202 124
rect 196 119 202 120
rect 127 110 129 113
rect 143 110 145 113
rect 153 110 155 113
rect 163 110 165 113
rect 116 108 129 110
rect 135 108 145 110
rect 149 109 155 110
rect 60 100 66 101
rect 119 100 121 108
rect 135 104 137 108
rect 149 105 150 109
rect 154 105 155 109
rect 149 104 155 105
rect 159 109 165 110
rect 159 105 160 109
rect 164 105 165 109
rect 200 110 202 119
rect 247 140 249 144
rect 227 131 229 135
rect 237 131 239 135
rect 456 142 458 146
rect 380 134 386 135
rect 283 132 289 133
rect 273 124 275 129
rect 283 128 284 132
rect 288 128 289 132
rect 283 127 289 128
rect 211 110 213 113
rect 227 110 229 113
rect 237 110 239 113
rect 247 110 249 113
rect 283 122 285 127
rect 293 122 295 127
rect 370 126 372 131
rect 380 130 381 134
rect 385 130 386 134
rect 380 129 386 130
rect 380 124 382 129
rect 390 124 392 129
rect 441 126 447 127
rect 441 122 442 126
rect 446 122 447 126
rect 441 121 447 122
rect 200 108 213 110
rect 219 108 229 110
rect 233 109 239 110
rect 159 104 165 105
rect 128 103 137 104
rect 60 96 61 100
rect 65 96 66 100
rect 60 95 66 96
rect 60 92 62 95
rect 41 85 43 89
rect 128 99 129 103
rect 133 99 137 103
rect 153 100 155 104
rect 128 98 137 99
rect 135 95 137 98
rect 145 95 147 100
rect 153 98 157 100
rect 155 95 157 98
rect 162 95 164 104
rect 203 100 205 108
rect 219 104 221 108
rect 233 105 234 109
rect 238 105 239 109
rect 233 104 239 105
rect 243 109 249 110
rect 243 105 244 109
rect 248 105 249 109
rect 243 104 249 105
rect 273 109 275 112
rect 283 109 285 112
rect 273 108 279 109
rect 273 104 274 108
rect 278 104 279 108
rect 283 106 287 109
rect 212 103 221 104
rect 119 88 121 91
rect 119 86 124 88
rect 53 78 55 83
rect 60 78 62 83
rect 122 78 124 86
rect 135 82 137 86
rect 145 78 147 86
rect 212 99 213 103
rect 217 99 221 103
rect 237 100 239 104
rect 212 98 221 99
rect 219 95 221 98
rect 229 95 231 100
rect 237 98 241 100
rect 239 95 241 98
rect 246 95 248 104
rect 273 103 279 104
rect 273 95 275 103
rect 203 88 205 91
rect 203 86 208 88
rect 155 78 157 83
rect 162 78 164 83
rect 122 76 147 78
rect 206 78 208 86
rect 219 82 221 86
rect 229 78 231 86
rect 285 92 287 106
rect 293 101 295 112
rect 370 111 372 114
rect 380 111 382 114
rect 370 110 376 111
rect 370 106 371 110
rect 375 106 376 110
rect 380 108 384 111
rect 370 105 376 106
rect 292 100 298 101
rect 292 96 293 100
rect 297 96 298 100
rect 370 97 372 105
rect 292 95 298 96
rect 292 92 294 95
rect 273 85 275 89
rect 382 94 384 108
rect 390 103 392 114
rect 445 112 447 121
rect 492 142 494 146
rect 540 142 542 146
rect 472 133 474 137
rect 482 133 484 137
rect 525 126 531 127
rect 525 122 526 126
rect 530 122 531 126
rect 525 121 531 122
rect 456 112 458 115
rect 472 112 474 115
rect 482 112 484 115
rect 492 112 494 115
rect 445 110 458 112
rect 464 110 474 112
rect 478 111 484 112
rect 389 102 395 103
rect 448 102 450 110
rect 464 106 466 110
rect 478 107 479 111
rect 483 107 484 111
rect 478 106 484 107
rect 488 111 494 112
rect 488 107 489 111
rect 493 107 494 111
rect 529 112 531 121
rect 576 142 578 146
rect 556 133 558 137
rect 566 133 568 137
rect 783 145 785 149
rect 707 137 713 138
rect 612 134 618 135
rect 602 126 604 131
rect 612 130 613 134
rect 617 130 618 134
rect 612 129 618 130
rect 697 129 699 134
rect 707 133 708 137
rect 712 133 713 137
rect 707 132 713 133
rect 540 112 542 115
rect 556 112 558 115
rect 566 112 568 115
rect 576 112 578 115
rect 612 124 614 129
rect 622 124 624 129
rect 707 127 709 132
rect 717 127 719 132
rect 768 129 774 130
rect 768 125 769 129
rect 773 125 774 129
rect 768 124 774 125
rect 697 114 699 117
rect 707 114 709 117
rect 529 110 542 112
rect 548 110 558 112
rect 562 111 568 112
rect 488 106 494 107
rect 457 105 466 106
rect 389 98 390 102
rect 394 98 395 102
rect 389 97 395 98
rect 389 94 391 97
rect 370 87 372 91
rect 457 101 458 105
rect 462 101 466 105
rect 482 102 484 106
rect 457 100 466 101
rect 464 97 466 100
rect 474 97 476 102
rect 482 100 486 102
rect 484 97 486 100
rect 491 97 493 106
rect 532 102 534 110
rect 548 106 550 110
rect 562 107 563 111
rect 567 107 568 111
rect 562 106 568 107
rect 572 111 578 112
rect 572 107 573 111
rect 577 107 578 111
rect 572 106 578 107
rect 602 111 604 114
rect 612 111 614 114
rect 602 110 608 111
rect 602 106 603 110
rect 607 106 608 110
rect 612 108 616 111
rect 541 105 550 106
rect 448 90 450 93
rect 448 88 453 90
rect 239 78 241 83
rect 246 78 248 83
rect 206 76 231 78
rect 285 78 287 83
rect 292 78 294 83
rect 382 80 384 85
rect 389 80 391 85
rect 451 80 453 88
rect 464 84 466 88
rect 474 80 476 88
rect 541 101 542 105
rect 546 101 550 105
rect 566 102 568 106
rect 541 100 550 101
rect 548 97 550 100
rect 558 97 560 102
rect 566 100 570 102
rect 568 97 570 100
rect 575 97 577 106
rect 602 105 608 106
rect 602 97 604 105
rect 532 90 534 93
rect 532 88 537 90
rect 484 80 486 85
rect 491 80 493 85
rect 451 78 476 80
rect 535 80 537 88
rect 548 84 550 88
rect 558 80 560 88
rect 614 94 616 108
rect 622 103 624 114
rect 697 113 703 114
rect 697 109 698 113
rect 702 109 703 113
rect 707 111 711 114
rect 697 108 703 109
rect 621 102 627 103
rect 621 98 622 102
rect 626 98 627 102
rect 697 100 699 108
rect 621 97 627 98
rect 621 94 623 97
rect 709 97 711 111
rect 717 106 719 117
rect 772 115 774 124
rect 819 145 821 149
rect 867 145 869 149
rect 799 136 801 140
rect 809 136 811 140
rect 852 129 858 130
rect 852 125 853 129
rect 857 125 858 129
rect 852 124 858 125
rect 783 115 785 118
rect 799 115 801 118
rect 809 115 811 118
rect 819 115 821 118
rect 772 113 785 115
rect 791 113 801 115
rect 805 114 811 115
rect 716 105 722 106
rect 775 105 777 113
rect 791 109 793 113
rect 805 110 806 114
rect 810 110 811 114
rect 805 109 811 110
rect 815 114 821 115
rect 815 110 816 114
rect 820 110 821 114
rect 856 115 858 124
rect 903 145 905 149
rect 883 136 885 140
rect 893 136 895 140
rect 939 137 945 138
rect 929 129 931 134
rect 939 133 940 137
rect 944 133 945 137
rect 939 132 945 133
rect 867 115 869 118
rect 883 115 885 118
rect 893 115 895 118
rect 903 115 905 118
rect 939 127 941 132
rect 949 127 951 132
rect 856 113 869 115
rect 875 113 885 115
rect 889 114 895 115
rect 815 109 821 110
rect 784 108 793 109
rect 716 101 717 105
rect 721 101 722 105
rect 716 100 722 101
rect 716 97 718 100
rect 602 87 604 91
rect 697 90 699 94
rect 784 104 785 108
rect 789 104 793 108
rect 809 105 811 109
rect 784 103 793 104
rect 791 100 793 103
rect 801 100 803 105
rect 809 103 813 105
rect 811 100 813 103
rect 818 100 820 109
rect 859 105 861 113
rect 875 109 877 113
rect 889 110 890 114
rect 894 110 895 114
rect 889 109 895 110
rect 899 114 905 115
rect 899 110 900 114
rect 904 110 905 114
rect 899 109 905 110
rect 929 114 931 117
rect 939 114 941 117
rect 929 113 935 114
rect 929 109 930 113
rect 934 109 935 113
rect 939 111 943 114
rect 868 108 877 109
rect 775 93 777 96
rect 775 91 780 93
rect 568 80 570 85
rect 575 80 577 85
rect 535 78 560 80
rect 614 80 616 85
rect 621 80 623 85
rect 709 83 711 88
rect 716 83 718 88
rect 778 83 780 91
rect 791 87 793 91
rect 801 83 803 91
rect 868 104 869 108
rect 873 104 877 108
rect 893 105 895 109
rect 868 103 877 104
rect 875 100 877 103
rect 885 100 887 105
rect 893 103 897 105
rect 895 100 897 103
rect 902 100 904 109
rect 929 108 935 109
rect 929 100 931 108
rect 859 93 861 96
rect 859 91 864 93
rect 811 83 813 88
rect 818 83 820 88
rect 778 81 803 83
rect 862 83 864 91
rect 875 87 877 91
rect 885 83 887 91
rect 941 97 943 111
rect 949 106 951 117
rect 948 105 954 106
rect 948 101 949 105
rect 953 101 954 105
rect 948 100 954 101
rect 948 97 950 100
rect 929 90 931 94
rect 895 83 897 88
rect 902 83 904 88
rect 862 81 887 83
rect 941 83 943 88
rect 948 83 950 88
rect 134 61 136 65
rect 144 61 146 65
rect 154 61 156 65
rect 463 63 465 67
rect 473 63 475 67
rect 483 63 485 67
rect 790 66 792 70
rect 800 66 802 70
rect 810 66 812 70
rect 134 47 136 55
rect 130 46 136 47
rect 144 46 146 55
rect 154 46 156 55
rect 463 49 465 57
rect 130 42 131 46
rect 135 42 136 46
rect 150 45 156 46
rect 130 41 136 42
rect 134 28 136 41
rect 144 39 146 42
rect 150 41 151 45
rect 155 41 156 45
rect 459 48 465 49
rect 473 48 475 57
rect 483 48 485 57
rect 790 52 792 60
rect 459 44 460 48
rect 464 44 465 48
rect 479 47 485 48
rect 459 43 465 44
rect 150 40 156 41
rect 140 38 146 39
rect 140 34 141 38
rect 145 34 146 38
rect 140 33 146 34
rect 141 28 143 33
rect 154 31 156 40
rect 463 30 465 43
rect 473 41 475 44
rect 479 43 480 47
rect 484 43 485 47
rect 786 51 792 52
rect 800 51 802 60
rect 810 51 812 60
rect 786 47 787 51
rect 791 47 792 51
rect 806 50 812 51
rect 786 46 792 47
rect 479 42 485 43
rect 469 40 475 41
rect 469 36 470 40
rect 474 36 475 40
rect 469 35 475 36
rect 470 30 472 35
rect 483 33 485 42
rect 790 33 792 46
rect 800 44 802 47
rect 806 46 807 50
rect 811 46 812 50
rect 806 45 812 46
rect 796 43 802 44
rect 796 39 797 43
rect 801 39 802 43
rect 796 38 802 39
rect 797 33 799 38
rect 810 36 812 45
rect 154 15 156 19
rect 483 17 485 21
rect 810 20 812 24
rect 134 6 136 10
rect 141 6 143 10
rect 463 8 465 12
rect 470 8 472 12
rect 790 11 792 15
rect 797 11 799 15
rect 126 -6 128 -2
rect 50 -14 56 -13
rect 40 -22 42 -17
rect 50 -18 51 -14
rect 55 -18 56 -14
rect 50 -19 56 -18
rect 50 -24 52 -19
rect 60 -24 62 -19
rect 111 -22 117 -21
rect 111 -26 112 -22
rect 116 -26 117 -22
rect 111 -27 117 -26
rect 40 -37 42 -34
rect 50 -37 52 -34
rect 40 -38 46 -37
rect 40 -42 41 -38
rect 45 -42 46 -38
rect 50 -40 54 -37
rect 40 -43 46 -42
rect 40 -51 42 -43
rect 52 -54 54 -40
rect 60 -45 62 -34
rect 115 -36 117 -27
rect 162 -6 164 -2
rect 210 -6 212 -2
rect 142 -15 144 -11
rect 152 -15 154 -11
rect 195 -22 201 -21
rect 195 -26 196 -22
rect 200 -26 201 -22
rect 195 -27 201 -26
rect 126 -36 128 -33
rect 142 -36 144 -33
rect 152 -36 154 -33
rect 162 -36 164 -33
rect 115 -38 128 -36
rect 134 -38 144 -36
rect 148 -37 154 -36
rect 59 -46 65 -45
rect 118 -46 120 -38
rect 134 -42 136 -38
rect 148 -41 149 -37
rect 153 -41 154 -37
rect 148 -42 154 -41
rect 158 -37 164 -36
rect 158 -41 159 -37
rect 163 -41 164 -37
rect 199 -36 201 -27
rect 246 -6 248 -2
rect 226 -15 228 -11
rect 236 -15 238 -11
rect 455 -4 457 0
rect 379 -12 385 -11
rect 282 -14 288 -13
rect 272 -22 274 -17
rect 282 -18 283 -14
rect 287 -18 288 -14
rect 282 -19 288 -18
rect 210 -36 212 -33
rect 226 -36 228 -33
rect 236 -36 238 -33
rect 246 -36 248 -33
rect 282 -24 284 -19
rect 292 -24 294 -19
rect 369 -20 371 -15
rect 379 -16 380 -12
rect 384 -16 385 -12
rect 379 -17 385 -16
rect 379 -22 381 -17
rect 389 -22 391 -17
rect 440 -20 446 -19
rect 440 -24 441 -20
rect 445 -24 446 -20
rect 440 -25 446 -24
rect 199 -38 212 -36
rect 218 -38 228 -36
rect 232 -37 238 -36
rect 158 -42 164 -41
rect 127 -43 136 -42
rect 59 -50 60 -46
rect 64 -50 65 -46
rect 59 -51 65 -50
rect 59 -54 61 -51
rect 40 -61 42 -57
rect 127 -47 128 -43
rect 132 -47 136 -43
rect 152 -46 154 -42
rect 127 -48 136 -47
rect 134 -51 136 -48
rect 144 -51 146 -46
rect 152 -48 156 -46
rect 154 -51 156 -48
rect 161 -51 163 -42
rect 202 -46 204 -38
rect 218 -42 220 -38
rect 232 -41 233 -37
rect 237 -41 238 -37
rect 232 -42 238 -41
rect 242 -37 248 -36
rect 242 -41 243 -37
rect 247 -41 248 -37
rect 242 -42 248 -41
rect 272 -37 274 -34
rect 282 -37 284 -34
rect 272 -38 278 -37
rect 272 -42 273 -38
rect 277 -42 278 -38
rect 282 -40 286 -37
rect 211 -43 220 -42
rect 118 -58 120 -55
rect 118 -60 123 -58
rect 52 -68 54 -63
rect 59 -68 61 -63
rect 121 -68 123 -60
rect 134 -64 136 -60
rect 144 -68 146 -60
rect 211 -47 212 -43
rect 216 -47 220 -43
rect 236 -46 238 -42
rect 211 -48 220 -47
rect 218 -51 220 -48
rect 228 -51 230 -46
rect 236 -48 240 -46
rect 238 -51 240 -48
rect 245 -51 247 -42
rect 272 -43 278 -42
rect 272 -51 274 -43
rect 202 -58 204 -55
rect 202 -60 207 -58
rect 154 -68 156 -63
rect 161 -68 163 -63
rect 121 -70 146 -68
rect 205 -68 207 -60
rect 218 -64 220 -60
rect 228 -68 230 -60
rect 284 -54 286 -40
rect 292 -45 294 -34
rect 369 -35 371 -32
rect 379 -35 381 -32
rect 369 -36 375 -35
rect 369 -40 370 -36
rect 374 -40 375 -36
rect 379 -38 383 -35
rect 369 -41 375 -40
rect 291 -46 297 -45
rect 291 -50 292 -46
rect 296 -50 297 -46
rect 369 -49 371 -41
rect 291 -51 297 -50
rect 291 -54 293 -51
rect 272 -61 274 -57
rect 381 -52 383 -38
rect 389 -43 391 -32
rect 444 -34 446 -25
rect 491 -4 493 0
rect 539 -4 541 0
rect 471 -13 473 -9
rect 481 -13 483 -9
rect 524 -20 530 -19
rect 524 -24 525 -20
rect 529 -24 530 -20
rect 524 -25 530 -24
rect 455 -34 457 -31
rect 471 -34 473 -31
rect 481 -34 483 -31
rect 491 -34 493 -31
rect 444 -36 457 -34
rect 463 -36 473 -34
rect 477 -35 483 -34
rect 388 -44 394 -43
rect 447 -44 449 -36
rect 463 -40 465 -36
rect 477 -39 478 -35
rect 482 -39 483 -35
rect 477 -40 483 -39
rect 487 -35 493 -34
rect 487 -39 488 -35
rect 492 -39 493 -35
rect 528 -34 530 -25
rect 575 -4 577 0
rect 555 -13 557 -9
rect 565 -13 567 -9
rect 782 -1 784 3
rect 706 -9 712 -8
rect 611 -12 617 -11
rect 601 -20 603 -15
rect 611 -16 612 -12
rect 616 -16 617 -12
rect 611 -17 617 -16
rect 696 -17 698 -12
rect 706 -13 707 -9
rect 711 -13 712 -9
rect 706 -14 712 -13
rect 539 -34 541 -31
rect 555 -34 557 -31
rect 565 -34 567 -31
rect 575 -34 577 -31
rect 611 -22 613 -17
rect 621 -22 623 -17
rect 706 -19 708 -14
rect 716 -19 718 -14
rect 767 -17 773 -16
rect 767 -21 768 -17
rect 772 -21 773 -17
rect 767 -22 773 -21
rect 696 -32 698 -29
rect 706 -32 708 -29
rect 528 -36 541 -34
rect 547 -36 557 -34
rect 561 -35 567 -34
rect 487 -40 493 -39
rect 456 -41 465 -40
rect 388 -48 389 -44
rect 393 -48 394 -44
rect 388 -49 394 -48
rect 388 -52 390 -49
rect 369 -59 371 -55
rect 456 -45 457 -41
rect 461 -45 465 -41
rect 481 -44 483 -40
rect 456 -46 465 -45
rect 463 -49 465 -46
rect 473 -49 475 -44
rect 481 -46 485 -44
rect 483 -49 485 -46
rect 490 -49 492 -40
rect 531 -44 533 -36
rect 547 -40 549 -36
rect 561 -39 562 -35
rect 566 -39 567 -35
rect 561 -40 567 -39
rect 571 -35 577 -34
rect 571 -39 572 -35
rect 576 -39 577 -35
rect 571 -40 577 -39
rect 601 -35 603 -32
rect 611 -35 613 -32
rect 601 -36 607 -35
rect 601 -40 602 -36
rect 606 -40 607 -36
rect 611 -38 615 -35
rect 540 -41 549 -40
rect 447 -56 449 -53
rect 447 -58 452 -56
rect 238 -68 240 -63
rect 245 -68 247 -63
rect 205 -70 230 -68
rect 284 -68 286 -63
rect 291 -68 293 -63
rect 381 -66 383 -61
rect 388 -66 390 -61
rect 450 -66 452 -58
rect 463 -62 465 -58
rect 473 -66 475 -58
rect 540 -45 541 -41
rect 545 -45 549 -41
rect 565 -44 567 -40
rect 540 -46 549 -45
rect 547 -49 549 -46
rect 557 -49 559 -44
rect 565 -46 569 -44
rect 567 -49 569 -46
rect 574 -49 576 -40
rect 601 -41 607 -40
rect 601 -49 603 -41
rect 531 -56 533 -53
rect 531 -58 536 -56
rect 483 -66 485 -61
rect 490 -66 492 -61
rect 450 -68 475 -66
rect 534 -66 536 -58
rect 547 -62 549 -58
rect 557 -66 559 -58
rect 613 -52 615 -38
rect 621 -43 623 -32
rect 696 -33 702 -32
rect 696 -37 697 -33
rect 701 -37 702 -33
rect 706 -35 710 -32
rect 696 -38 702 -37
rect 620 -44 626 -43
rect 620 -48 621 -44
rect 625 -48 626 -44
rect 696 -46 698 -38
rect 620 -49 626 -48
rect 620 -52 622 -49
rect 708 -49 710 -35
rect 716 -40 718 -29
rect 771 -31 773 -22
rect 818 -1 820 3
rect 866 -1 868 3
rect 798 -10 800 -6
rect 808 -10 810 -6
rect 851 -17 857 -16
rect 851 -21 852 -17
rect 856 -21 857 -17
rect 851 -22 857 -21
rect 782 -31 784 -28
rect 798 -31 800 -28
rect 808 -31 810 -28
rect 818 -31 820 -28
rect 771 -33 784 -31
rect 790 -33 800 -31
rect 804 -32 810 -31
rect 715 -41 721 -40
rect 774 -41 776 -33
rect 790 -37 792 -33
rect 804 -36 805 -32
rect 809 -36 810 -32
rect 804 -37 810 -36
rect 814 -32 820 -31
rect 814 -36 815 -32
rect 819 -36 820 -32
rect 855 -31 857 -22
rect 902 -1 904 3
rect 882 -10 884 -6
rect 892 -10 894 -6
rect 938 -9 944 -8
rect 928 -17 930 -12
rect 938 -13 939 -9
rect 943 -13 944 -9
rect 938 -14 944 -13
rect 866 -31 868 -28
rect 882 -31 884 -28
rect 892 -31 894 -28
rect 902 -31 904 -28
rect 938 -19 940 -14
rect 948 -19 950 -14
rect 855 -33 868 -31
rect 874 -33 884 -31
rect 888 -32 894 -31
rect 814 -37 820 -36
rect 783 -38 792 -37
rect 715 -45 716 -41
rect 720 -45 721 -41
rect 715 -46 721 -45
rect 715 -49 717 -46
rect 601 -59 603 -55
rect 696 -56 698 -52
rect 783 -42 784 -38
rect 788 -42 792 -38
rect 808 -41 810 -37
rect 783 -43 792 -42
rect 790 -46 792 -43
rect 800 -46 802 -41
rect 808 -43 812 -41
rect 810 -46 812 -43
rect 817 -46 819 -37
rect 858 -41 860 -33
rect 874 -37 876 -33
rect 888 -36 889 -32
rect 893 -36 894 -32
rect 888 -37 894 -36
rect 898 -32 904 -31
rect 898 -36 899 -32
rect 903 -36 904 -32
rect 898 -37 904 -36
rect 928 -32 930 -29
rect 938 -32 940 -29
rect 928 -33 934 -32
rect 928 -37 929 -33
rect 933 -37 934 -33
rect 938 -35 942 -32
rect 867 -38 876 -37
rect 774 -53 776 -50
rect 774 -55 779 -53
rect 567 -66 569 -61
rect 574 -66 576 -61
rect 534 -68 559 -66
rect 613 -66 615 -61
rect 620 -66 622 -61
rect 708 -63 710 -58
rect 715 -63 717 -58
rect 777 -63 779 -55
rect 790 -59 792 -55
rect 800 -63 802 -55
rect 867 -42 868 -38
rect 872 -42 876 -38
rect 892 -41 894 -37
rect 867 -43 876 -42
rect 874 -46 876 -43
rect 884 -46 886 -41
rect 892 -43 896 -41
rect 894 -46 896 -43
rect 901 -46 903 -37
rect 928 -38 934 -37
rect 928 -46 930 -38
rect 858 -53 860 -50
rect 858 -55 863 -53
rect 810 -63 812 -58
rect 817 -63 819 -58
rect 777 -65 802 -63
rect 861 -63 863 -55
rect 874 -59 876 -55
rect 884 -63 886 -55
rect 940 -49 942 -35
rect 948 -40 950 -29
rect 947 -41 953 -40
rect 947 -45 948 -41
rect 952 -45 953 -41
rect 947 -46 953 -45
rect 947 -49 949 -46
rect 928 -56 930 -52
rect 894 -63 896 -58
rect 901 -63 903 -58
rect 861 -65 886 -63
rect 940 -63 942 -58
rect 947 -63 949 -58
rect 133 -85 135 -81
rect 143 -85 145 -81
rect 153 -85 155 -81
rect 462 -83 464 -79
rect 472 -83 474 -79
rect 482 -83 484 -79
rect 789 -80 791 -76
rect 799 -80 801 -76
rect 809 -80 811 -76
rect 133 -99 135 -91
rect 129 -100 135 -99
rect 143 -100 145 -91
rect 153 -100 155 -91
rect 462 -97 464 -89
rect 129 -104 130 -100
rect 134 -104 135 -100
rect 149 -101 155 -100
rect 129 -105 135 -104
rect 133 -118 135 -105
rect 143 -107 145 -104
rect 149 -105 150 -101
rect 154 -105 155 -101
rect 458 -98 464 -97
rect 472 -98 474 -89
rect 482 -98 484 -89
rect 789 -94 791 -86
rect 458 -102 459 -98
rect 463 -102 464 -98
rect 478 -99 484 -98
rect 458 -103 464 -102
rect 149 -106 155 -105
rect 139 -108 145 -107
rect 139 -112 140 -108
rect 144 -112 145 -108
rect 139 -113 145 -112
rect 140 -118 142 -113
rect 153 -115 155 -106
rect 462 -116 464 -103
rect 472 -105 474 -102
rect 478 -103 479 -99
rect 483 -103 484 -99
rect 785 -95 791 -94
rect 799 -95 801 -86
rect 809 -95 811 -86
rect 785 -99 786 -95
rect 790 -99 791 -95
rect 805 -96 811 -95
rect 785 -100 791 -99
rect 478 -104 484 -103
rect 468 -106 474 -105
rect 468 -110 469 -106
rect 473 -110 474 -106
rect 468 -111 474 -110
rect 469 -116 471 -111
rect 482 -113 484 -104
rect 789 -113 791 -100
rect 799 -102 801 -99
rect 805 -100 806 -96
rect 810 -100 811 -96
rect 805 -101 811 -100
rect 795 -103 801 -102
rect 795 -107 796 -103
rect 800 -107 801 -103
rect 795 -108 801 -107
rect 796 -113 798 -108
rect 809 -110 811 -101
rect 153 -131 155 -127
rect 482 -129 484 -125
rect 809 -126 811 -122
rect 133 -140 135 -136
rect 140 -140 142 -136
rect 462 -138 464 -134
rect 469 -138 471 -134
rect 789 -135 791 -131
rect 796 -135 798 -131
rect 334 -163 336 -159
rect 344 -161 346 -156
rect 354 -161 356 -156
rect 427 -163 429 -159
rect 437 -161 439 -156
rect 447 -161 449 -156
rect 334 -185 336 -181
rect 344 -185 346 -174
rect 354 -177 356 -174
rect 354 -178 360 -177
rect 354 -182 355 -178
rect 359 -182 360 -178
rect 514 -163 516 -159
rect 524 -161 526 -156
rect 534 -161 536 -156
rect 354 -183 360 -182
rect 334 -186 340 -185
rect 334 -190 335 -186
rect 339 -190 340 -186
rect 334 -191 340 -190
rect 344 -186 350 -185
rect 344 -190 345 -186
rect 349 -190 350 -186
rect 344 -191 350 -190
rect 334 -196 336 -191
rect 347 -196 349 -191
rect 354 -196 356 -183
rect 427 -185 429 -181
rect 437 -185 439 -174
rect 447 -177 449 -174
rect 447 -178 453 -177
rect 447 -182 448 -178
rect 452 -182 453 -178
rect 447 -183 453 -182
rect 427 -186 433 -185
rect 427 -190 428 -186
rect 432 -190 433 -186
rect 427 -191 433 -190
rect 437 -186 443 -185
rect 437 -190 438 -186
rect 442 -190 443 -186
rect 437 -191 443 -190
rect 427 -196 429 -191
rect 440 -196 442 -191
rect 447 -196 449 -183
rect 514 -185 516 -181
rect 524 -185 526 -174
rect 534 -177 536 -174
rect 534 -178 540 -177
rect 534 -182 535 -178
rect 539 -182 540 -178
rect 534 -183 540 -182
rect 514 -186 520 -185
rect 514 -190 515 -186
rect 519 -190 520 -186
rect 514 -191 520 -190
rect 524 -186 530 -185
rect 524 -190 525 -186
rect 529 -190 530 -186
rect 524 -191 530 -190
rect 514 -196 516 -191
rect 527 -196 529 -191
rect 534 -196 536 -183
rect 334 -209 336 -205
rect 347 -212 349 -207
rect 354 -212 356 -207
rect 427 -209 429 -205
rect 440 -212 442 -207
rect 447 -212 449 -207
rect 514 -209 516 -205
rect 527 -212 529 -207
rect 534 -212 536 -207
<< ndiffusion >>
rect 130 221 137 222
rect 130 217 132 221
rect 136 217 137 221
rect 130 212 137 217
rect 217 221 224 222
rect 217 217 219 221
rect 223 217 224 221
rect 112 211 119 212
rect 112 207 113 211
rect 117 207 119 211
rect 112 206 119 207
rect 114 201 119 206
rect 121 201 126 212
rect 128 210 137 212
rect 217 212 224 217
rect 310 221 317 222
rect 310 217 312 221
rect 316 217 317 221
rect 199 211 206 212
rect 128 201 139 210
rect 141 209 148 210
rect 141 205 143 209
rect 147 205 148 209
rect 199 207 200 211
rect 204 207 206 211
rect 199 206 206 207
rect 141 204 148 205
rect 141 201 146 204
rect 201 201 206 206
rect 208 201 213 212
rect 215 210 224 212
rect 310 212 317 217
rect 543 223 550 224
rect 543 219 544 223
rect 548 219 550 223
rect 292 211 299 212
rect 215 201 226 210
rect 228 209 235 210
rect 228 205 230 209
rect 234 205 235 209
rect 292 207 293 211
rect 297 207 299 211
rect 292 206 299 207
rect 228 204 235 205
rect 228 201 233 204
rect 294 201 299 206
rect 301 201 306 212
rect 308 210 317 212
rect 543 214 550 219
rect 636 223 643 224
rect 636 219 637 223
rect 641 219 643 223
rect 543 212 552 214
rect 532 211 539 212
rect 308 201 319 210
rect 321 209 328 210
rect 321 205 323 209
rect 327 205 328 209
rect 532 207 533 211
rect 537 207 539 211
rect 532 206 539 207
rect 321 204 328 205
rect 321 201 326 204
rect 534 203 539 206
rect 541 203 552 212
rect 554 203 559 214
rect 561 213 568 214
rect 561 209 563 213
rect 567 209 568 213
rect 636 214 643 219
rect 723 223 730 224
rect 723 219 724 223
rect 728 219 730 223
rect 636 212 645 214
rect 561 208 568 209
rect 625 211 632 212
rect 561 203 566 208
rect 625 207 626 211
rect 630 207 632 211
rect 625 206 632 207
rect 627 203 632 206
rect 634 203 645 212
rect 647 203 652 214
rect 654 213 661 214
rect 654 209 656 213
rect 660 209 661 213
rect 723 214 730 219
rect 723 212 732 214
rect 654 208 661 209
rect 712 211 719 212
rect 654 203 659 208
rect 712 207 713 211
rect 717 207 719 211
rect 712 206 719 207
rect 714 203 719 206
rect 721 203 732 212
rect 734 203 739 214
rect 741 213 748 214
rect 741 209 743 213
rect 747 209 748 213
rect 741 208 748 209
rect 741 203 746 208
rect 34 94 41 95
rect 34 90 35 94
rect 39 90 41 94
rect 34 89 41 90
rect 43 92 51 95
rect 112 99 119 100
rect 112 95 113 99
rect 117 95 119 99
rect 112 94 119 95
rect 43 89 53 92
rect 45 83 53 89
rect 55 83 60 92
rect 62 91 69 92
rect 114 91 119 94
rect 121 95 126 100
rect 196 99 203 100
rect 196 95 197 99
rect 201 95 203 99
rect 121 91 135 95
rect 62 87 64 91
rect 68 87 69 91
rect 62 86 69 87
rect 126 87 127 91
rect 131 87 135 91
rect 126 86 135 87
rect 137 94 145 95
rect 137 90 139 94
rect 143 90 145 94
rect 137 86 145 90
rect 147 92 155 95
rect 147 88 149 92
rect 153 88 155 92
rect 147 86 155 88
rect 62 83 67 86
rect 45 82 51 83
rect 45 78 46 82
rect 50 78 51 82
rect 45 77 51 78
rect 150 83 155 86
rect 157 83 162 95
rect 164 83 172 95
rect 196 94 203 95
rect 198 91 203 94
rect 205 95 210 100
rect 205 91 219 95
rect 210 87 211 91
rect 215 87 219 91
rect 210 86 219 87
rect 221 94 229 95
rect 221 90 223 94
rect 227 90 229 94
rect 221 86 229 90
rect 231 92 239 95
rect 231 88 233 92
rect 237 88 239 92
rect 231 86 239 88
rect 166 82 172 83
rect 166 78 167 82
rect 171 78 172 82
rect 166 77 172 78
rect 234 83 239 86
rect 241 83 246 95
rect 248 83 256 95
rect 266 94 273 95
rect 266 90 267 94
rect 271 90 273 94
rect 266 89 273 90
rect 275 92 283 95
rect 363 96 370 97
rect 363 92 364 96
rect 368 92 370 96
rect 275 89 285 92
rect 277 83 285 89
rect 287 83 292 92
rect 294 91 301 92
rect 363 91 370 92
rect 372 94 380 97
rect 441 101 448 102
rect 441 97 442 101
rect 446 97 448 101
rect 441 96 448 97
rect 372 91 382 94
rect 294 87 296 91
rect 300 87 301 91
rect 294 86 301 87
rect 294 83 299 86
rect 374 85 382 91
rect 384 85 389 94
rect 391 93 398 94
rect 443 93 448 96
rect 450 97 455 102
rect 525 101 532 102
rect 525 97 526 101
rect 530 97 532 101
rect 450 93 464 97
rect 391 89 393 93
rect 397 89 398 93
rect 391 88 398 89
rect 455 89 456 93
rect 460 89 464 93
rect 455 88 464 89
rect 466 96 474 97
rect 466 92 468 96
rect 472 92 474 96
rect 466 88 474 92
rect 476 94 484 97
rect 476 90 478 94
rect 482 90 484 94
rect 476 88 484 90
rect 391 85 396 88
rect 250 82 256 83
rect 250 78 251 82
rect 255 78 256 82
rect 250 77 256 78
rect 277 82 283 83
rect 277 78 278 82
rect 282 78 283 82
rect 374 84 380 85
rect 374 80 375 84
rect 379 80 380 84
rect 374 79 380 80
rect 479 85 484 88
rect 486 85 491 97
rect 493 85 501 97
rect 525 96 532 97
rect 527 93 532 96
rect 534 97 539 102
rect 534 93 548 97
rect 539 89 540 93
rect 544 89 548 93
rect 539 88 548 89
rect 550 96 558 97
rect 550 92 552 96
rect 556 92 558 96
rect 550 88 558 92
rect 560 94 568 97
rect 560 90 562 94
rect 566 90 568 94
rect 560 88 568 90
rect 495 84 501 85
rect 495 80 496 84
rect 500 80 501 84
rect 495 79 501 80
rect 563 85 568 88
rect 570 85 575 97
rect 577 85 585 97
rect 595 96 602 97
rect 595 92 596 96
rect 600 92 602 96
rect 595 91 602 92
rect 604 94 612 97
rect 690 99 697 100
rect 690 95 691 99
rect 695 95 697 99
rect 690 94 697 95
rect 699 97 707 100
rect 768 104 775 105
rect 768 100 769 104
rect 773 100 775 104
rect 768 99 775 100
rect 699 94 709 97
rect 604 91 614 94
rect 606 85 614 91
rect 616 85 621 94
rect 623 93 630 94
rect 623 89 625 93
rect 629 89 630 93
rect 623 88 630 89
rect 701 88 709 94
rect 711 88 716 97
rect 718 96 725 97
rect 770 96 775 99
rect 777 100 782 105
rect 852 104 859 105
rect 852 100 853 104
rect 857 100 859 104
rect 777 96 791 100
rect 718 92 720 96
rect 724 92 725 96
rect 718 91 725 92
rect 782 92 783 96
rect 787 92 791 96
rect 782 91 791 92
rect 793 99 801 100
rect 793 95 795 99
rect 799 95 801 99
rect 793 91 801 95
rect 803 97 811 100
rect 803 93 805 97
rect 809 93 811 97
rect 803 91 811 93
rect 718 88 723 91
rect 623 85 628 88
rect 579 84 585 85
rect 579 80 580 84
rect 584 80 585 84
rect 579 79 585 80
rect 606 84 612 85
rect 606 80 607 84
rect 611 80 612 84
rect 701 87 707 88
rect 701 83 702 87
rect 706 83 707 87
rect 701 82 707 83
rect 806 88 811 91
rect 813 88 818 100
rect 820 88 828 100
rect 852 99 859 100
rect 854 96 859 99
rect 861 100 866 105
rect 861 96 875 100
rect 866 92 867 96
rect 871 92 875 96
rect 866 91 875 92
rect 877 99 885 100
rect 877 95 879 99
rect 883 95 885 99
rect 877 91 885 95
rect 887 97 895 100
rect 887 93 889 97
rect 893 93 895 97
rect 887 91 895 93
rect 822 87 828 88
rect 822 83 823 87
rect 827 83 828 87
rect 822 82 828 83
rect 890 88 895 91
rect 897 88 902 100
rect 904 88 912 100
rect 922 99 929 100
rect 922 95 923 99
rect 927 95 929 99
rect 922 94 929 95
rect 931 97 939 100
rect 931 94 941 97
rect 933 88 941 94
rect 943 88 948 97
rect 950 96 957 97
rect 950 92 952 96
rect 956 92 957 96
rect 950 91 957 92
rect 950 88 955 91
rect 906 87 912 88
rect 906 83 907 87
rect 911 83 912 87
rect 906 82 912 83
rect 933 87 939 88
rect 933 83 934 87
rect 938 83 939 87
rect 933 82 939 83
rect 606 79 612 80
rect 277 77 283 78
rect 783 65 790 66
rect 456 62 463 63
rect 127 60 134 61
rect 127 56 128 60
rect 132 56 134 60
rect 127 55 134 56
rect 136 60 144 61
rect 136 56 138 60
rect 142 56 144 60
rect 136 55 144 56
rect 146 60 154 61
rect 146 56 148 60
rect 152 56 154 60
rect 146 55 154 56
rect 156 60 163 61
rect 156 56 158 60
rect 162 56 163 60
rect 456 58 457 62
rect 461 58 463 62
rect 456 57 463 58
rect 465 62 473 63
rect 465 58 467 62
rect 471 58 473 62
rect 465 57 473 58
rect 475 62 483 63
rect 475 58 477 62
rect 481 58 483 62
rect 475 57 483 58
rect 485 62 492 63
rect 485 58 487 62
rect 491 58 492 62
rect 783 61 784 65
rect 788 61 790 65
rect 783 60 790 61
rect 792 65 800 66
rect 792 61 794 65
rect 798 61 800 65
rect 792 60 800 61
rect 802 65 810 66
rect 802 61 804 65
rect 808 61 810 65
rect 802 60 810 61
rect 812 65 819 66
rect 812 61 814 65
rect 818 61 819 65
rect 812 60 819 61
rect 485 57 492 58
rect 156 55 163 56
rect 33 -52 40 -51
rect 33 -56 34 -52
rect 38 -56 40 -52
rect 33 -57 40 -56
rect 42 -54 50 -51
rect 111 -47 118 -46
rect 111 -51 112 -47
rect 116 -51 118 -47
rect 111 -52 118 -51
rect 42 -57 52 -54
rect 44 -63 52 -57
rect 54 -63 59 -54
rect 61 -55 68 -54
rect 113 -55 118 -52
rect 120 -51 125 -46
rect 195 -47 202 -46
rect 195 -51 196 -47
rect 200 -51 202 -47
rect 120 -55 134 -51
rect 61 -59 63 -55
rect 67 -59 68 -55
rect 61 -60 68 -59
rect 125 -59 126 -55
rect 130 -59 134 -55
rect 125 -60 134 -59
rect 136 -52 144 -51
rect 136 -56 138 -52
rect 142 -56 144 -52
rect 136 -60 144 -56
rect 146 -54 154 -51
rect 146 -58 148 -54
rect 152 -58 154 -54
rect 146 -60 154 -58
rect 61 -63 66 -60
rect 44 -64 50 -63
rect 44 -68 45 -64
rect 49 -68 50 -64
rect 44 -69 50 -68
rect 149 -63 154 -60
rect 156 -63 161 -51
rect 163 -63 171 -51
rect 195 -52 202 -51
rect 197 -55 202 -52
rect 204 -51 209 -46
rect 204 -55 218 -51
rect 209 -59 210 -55
rect 214 -59 218 -55
rect 209 -60 218 -59
rect 220 -52 228 -51
rect 220 -56 222 -52
rect 226 -56 228 -52
rect 220 -60 228 -56
rect 230 -54 238 -51
rect 230 -58 232 -54
rect 236 -58 238 -54
rect 230 -60 238 -58
rect 165 -64 171 -63
rect 165 -68 166 -64
rect 170 -68 171 -64
rect 165 -69 171 -68
rect 233 -63 238 -60
rect 240 -63 245 -51
rect 247 -63 255 -51
rect 265 -52 272 -51
rect 265 -56 266 -52
rect 270 -56 272 -52
rect 265 -57 272 -56
rect 274 -54 282 -51
rect 362 -50 369 -49
rect 362 -54 363 -50
rect 367 -54 369 -50
rect 274 -57 284 -54
rect 276 -63 284 -57
rect 286 -63 291 -54
rect 293 -55 300 -54
rect 362 -55 369 -54
rect 371 -52 379 -49
rect 440 -45 447 -44
rect 440 -49 441 -45
rect 445 -49 447 -45
rect 440 -50 447 -49
rect 371 -55 381 -52
rect 293 -59 295 -55
rect 299 -59 300 -55
rect 293 -60 300 -59
rect 293 -63 298 -60
rect 373 -61 381 -55
rect 383 -61 388 -52
rect 390 -53 397 -52
rect 442 -53 447 -50
rect 449 -49 454 -44
rect 524 -45 531 -44
rect 524 -49 525 -45
rect 529 -49 531 -45
rect 449 -53 463 -49
rect 390 -57 392 -53
rect 396 -57 397 -53
rect 390 -58 397 -57
rect 454 -57 455 -53
rect 459 -57 463 -53
rect 454 -58 463 -57
rect 465 -50 473 -49
rect 465 -54 467 -50
rect 471 -54 473 -50
rect 465 -58 473 -54
rect 475 -52 483 -49
rect 475 -56 477 -52
rect 481 -56 483 -52
rect 475 -58 483 -56
rect 390 -61 395 -58
rect 249 -64 255 -63
rect 249 -68 250 -64
rect 254 -68 255 -64
rect 249 -69 255 -68
rect 276 -64 282 -63
rect 276 -68 277 -64
rect 281 -68 282 -64
rect 373 -62 379 -61
rect 373 -66 374 -62
rect 378 -66 379 -62
rect 373 -67 379 -66
rect 478 -61 483 -58
rect 485 -61 490 -49
rect 492 -61 500 -49
rect 524 -50 531 -49
rect 526 -53 531 -50
rect 533 -49 538 -44
rect 533 -53 547 -49
rect 538 -57 539 -53
rect 543 -57 547 -53
rect 538 -58 547 -57
rect 549 -50 557 -49
rect 549 -54 551 -50
rect 555 -54 557 -50
rect 549 -58 557 -54
rect 559 -52 567 -49
rect 559 -56 561 -52
rect 565 -56 567 -52
rect 559 -58 567 -56
rect 494 -62 500 -61
rect 494 -66 495 -62
rect 499 -66 500 -62
rect 494 -67 500 -66
rect 562 -61 567 -58
rect 569 -61 574 -49
rect 576 -61 584 -49
rect 594 -50 601 -49
rect 594 -54 595 -50
rect 599 -54 601 -50
rect 594 -55 601 -54
rect 603 -52 611 -49
rect 689 -47 696 -46
rect 689 -51 690 -47
rect 694 -51 696 -47
rect 689 -52 696 -51
rect 698 -49 706 -46
rect 767 -42 774 -41
rect 767 -46 768 -42
rect 772 -46 774 -42
rect 767 -47 774 -46
rect 698 -52 708 -49
rect 603 -55 613 -52
rect 605 -61 613 -55
rect 615 -61 620 -52
rect 622 -53 629 -52
rect 622 -57 624 -53
rect 628 -57 629 -53
rect 622 -58 629 -57
rect 700 -58 708 -52
rect 710 -58 715 -49
rect 717 -50 724 -49
rect 769 -50 774 -47
rect 776 -46 781 -41
rect 851 -42 858 -41
rect 851 -46 852 -42
rect 856 -46 858 -42
rect 776 -50 790 -46
rect 717 -54 719 -50
rect 723 -54 724 -50
rect 717 -55 724 -54
rect 781 -54 782 -50
rect 786 -54 790 -50
rect 781 -55 790 -54
rect 792 -47 800 -46
rect 792 -51 794 -47
rect 798 -51 800 -47
rect 792 -55 800 -51
rect 802 -49 810 -46
rect 802 -53 804 -49
rect 808 -53 810 -49
rect 802 -55 810 -53
rect 717 -58 722 -55
rect 622 -61 627 -58
rect 578 -62 584 -61
rect 578 -66 579 -62
rect 583 -66 584 -62
rect 578 -67 584 -66
rect 605 -62 611 -61
rect 605 -66 606 -62
rect 610 -66 611 -62
rect 700 -59 706 -58
rect 700 -63 701 -59
rect 705 -63 706 -59
rect 700 -64 706 -63
rect 805 -58 810 -55
rect 812 -58 817 -46
rect 819 -58 827 -46
rect 851 -47 858 -46
rect 853 -50 858 -47
rect 860 -46 865 -41
rect 860 -50 874 -46
rect 865 -54 866 -50
rect 870 -54 874 -50
rect 865 -55 874 -54
rect 876 -47 884 -46
rect 876 -51 878 -47
rect 882 -51 884 -47
rect 876 -55 884 -51
rect 886 -49 894 -46
rect 886 -53 888 -49
rect 892 -53 894 -49
rect 886 -55 894 -53
rect 821 -59 827 -58
rect 821 -63 822 -59
rect 826 -63 827 -59
rect 821 -64 827 -63
rect 889 -58 894 -55
rect 896 -58 901 -46
rect 903 -58 911 -46
rect 921 -47 928 -46
rect 921 -51 922 -47
rect 926 -51 928 -47
rect 921 -52 928 -51
rect 930 -49 938 -46
rect 930 -52 940 -49
rect 932 -58 940 -52
rect 942 -58 947 -49
rect 949 -50 956 -49
rect 949 -54 951 -50
rect 955 -54 956 -50
rect 949 -55 956 -54
rect 949 -58 954 -55
rect 905 -59 911 -58
rect 905 -63 906 -59
rect 910 -63 911 -59
rect 905 -64 911 -63
rect 932 -59 938 -58
rect 932 -63 933 -59
rect 937 -63 938 -59
rect 932 -64 938 -63
rect 605 -67 611 -66
rect 276 -69 282 -68
rect 782 -81 789 -80
rect 455 -84 462 -83
rect 126 -86 133 -85
rect 126 -90 127 -86
rect 131 -90 133 -86
rect 126 -91 133 -90
rect 135 -86 143 -85
rect 135 -90 137 -86
rect 141 -90 143 -86
rect 135 -91 143 -90
rect 145 -86 153 -85
rect 145 -90 147 -86
rect 151 -90 153 -86
rect 145 -91 153 -90
rect 155 -86 162 -85
rect 155 -90 157 -86
rect 161 -90 162 -86
rect 455 -88 456 -84
rect 460 -88 462 -84
rect 455 -89 462 -88
rect 464 -84 472 -83
rect 464 -88 466 -84
rect 470 -88 472 -84
rect 464 -89 472 -88
rect 474 -84 482 -83
rect 474 -88 476 -84
rect 480 -88 482 -84
rect 474 -89 482 -88
rect 484 -84 491 -83
rect 484 -88 486 -84
rect 490 -88 491 -84
rect 782 -85 783 -81
rect 787 -85 789 -81
rect 782 -86 789 -85
rect 791 -81 799 -80
rect 791 -85 793 -81
rect 797 -85 799 -81
rect 791 -86 799 -85
rect 801 -81 809 -80
rect 801 -85 803 -81
rect 807 -85 809 -81
rect 801 -86 809 -85
rect 811 -81 818 -80
rect 811 -85 813 -81
rect 817 -85 818 -81
rect 811 -86 818 -85
rect 484 -89 491 -88
rect 155 -91 162 -90
rect 329 -199 334 -196
rect 327 -200 334 -199
rect 327 -204 328 -200
rect 332 -204 334 -200
rect 327 -205 334 -204
rect 336 -205 347 -196
rect 338 -207 347 -205
rect 349 -207 354 -196
rect 356 -201 361 -196
rect 422 -199 427 -196
rect 420 -200 427 -199
rect 356 -202 363 -201
rect 356 -206 358 -202
rect 362 -206 363 -202
rect 420 -204 421 -200
rect 425 -204 427 -200
rect 420 -205 427 -204
rect 429 -205 440 -196
rect 356 -207 363 -206
rect 338 -212 345 -207
rect 431 -207 440 -205
rect 442 -207 447 -196
rect 449 -201 454 -196
rect 509 -199 514 -196
rect 507 -200 514 -199
rect 449 -202 456 -201
rect 449 -206 451 -202
rect 455 -206 456 -202
rect 507 -204 508 -200
rect 512 -204 514 -200
rect 507 -205 514 -204
rect 516 -205 527 -196
rect 449 -207 456 -206
rect 338 -216 339 -212
rect 343 -216 345 -212
rect 338 -217 345 -216
rect 431 -212 438 -207
rect 518 -207 527 -205
rect 529 -207 534 -196
rect 536 -201 541 -196
rect 536 -202 543 -201
rect 536 -206 538 -202
rect 542 -206 543 -202
rect 536 -207 543 -206
rect 431 -216 432 -212
rect 436 -216 438 -212
rect 431 -217 438 -216
rect 518 -212 525 -207
rect 518 -216 519 -212
rect 523 -216 525 -212
rect 518 -217 525 -216
<< pdiffusion >>
rect 133 179 139 186
rect 112 171 119 179
rect 112 167 113 171
rect 117 167 119 171
rect 112 166 119 167
rect 121 178 129 179
rect 121 174 123 178
rect 127 174 129 178
rect 121 171 129 174
rect 121 167 123 171
rect 127 167 129 171
rect 121 166 129 167
rect 131 173 139 179
rect 131 169 133 173
rect 137 169 139 173
rect 131 168 139 169
rect 141 185 148 186
rect 141 181 143 185
rect 147 181 148 185
rect 141 178 148 181
rect 220 179 226 186
rect 141 174 143 178
rect 147 174 148 178
rect 141 173 148 174
rect 141 168 146 173
rect 199 171 206 179
rect 131 166 137 168
rect 199 167 200 171
rect 204 167 206 171
rect 199 166 206 167
rect 208 178 216 179
rect 208 174 210 178
rect 214 174 216 178
rect 208 171 216 174
rect 208 167 210 171
rect 214 167 216 171
rect 208 166 216 167
rect 218 173 226 179
rect 218 169 220 173
rect 224 169 226 173
rect 218 168 226 169
rect 228 185 235 186
rect 228 181 230 185
rect 234 181 235 185
rect 228 178 235 181
rect 532 187 539 188
rect 313 179 319 186
rect 228 174 230 178
rect 234 174 235 178
rect 228 173 235 174
rect 228 168 233 173
rect 292 171 299 179
rect 218 166 224 168
rect 292 167 293 171
rect 297 167 299 171
rect 292 166 299 167
rect 301 178 309 179
rect 301 174 303 178
rect 307 174 309 178
rect 301 171 309 174
rect 301 167 303 171
rect 307 167 309 171
rect 301 166 309 167
rect 311 173 319 179
rect 311 169 313 173
rect 317 169 319 173
rect 311 168 319 169
rect 321 185 328 186
rect 321 181 323 185
rect 327 181 328 185
rect 321 178 328 181
rect 321 174 323 178
rect 327 174 328 178
rect 532 183 533 187
rect 537 183 539 187
rect 532 180 539 183
rect 532 176 533 180
rect 537 176 539 180
rect 532 175 539 176
rect 321 173 328 174
rect 321 168 326 173
rect 534 170 539 175
rect 541 181 547 188
rect 625 187 632 188
rect 625 183 626 187
rect 630 183 632 187
rect 541 175 549 181
rect 541 171 543 175
rect 547 171 549 175
rect 541 170 549 171
rect 311 166 317 168
rect 543 168 549 170
rect 551 180 559 181
rect 551 176 553 180
rect 557 176 559 180
rect 551 173 559 176
rect 551 169 553 173
rect 557 169 559 173
rect 551 168 559 169
rect 561 173 568 181
rect 625 180 632 183
rect 625 176 626 180
rect 630 176 632 180
rect 625 175 632 176
rect 561 169 563 173
rect 567 169 568 173
rect 627 170 632 175
rect 634 181 640 188
rect 712 187 719 188
rect 712 183 713 187
rect 717 183 719 187
rect 634 175 642 181
rect 634 171 636 175
rect 640 171 642 175
rect 634 170 642 171
rect 561 168 568 169
rect 636 168 642 170
rect 644 180 652 181
rect 644 176 646 180
rect 650 176 652 180
rect 644 173 652 176
rect 644 169 646 173
rect 650 169 652 173
rect 644 168 652 169
rect 654 173 661 181
rect 712 180 719 183
rect 712 176 713 180
rect 717 176 719 180
rect 712 175 719 176
rect 654 169 656 173
rect 660 169 661 173
rect 714 170 719 175
rect 721 181 727 188
rect 721 175 729 181
rect 721 171 723 175
rect 727 171 729 175
rect 721 170 729 171
rect 654 168 661 169
rect 723 168 729 170
rect 731 180 739 181
rect 731 176 733 180
rect 737 176 739 180
rect 731 173 739 176
rect 731 169 733 173
rect 737 169 739 173
rect 731 168 739 169
rect 741 173 748 181
rect 741 169 743 173
rect 747 169 748 173
rect 741 168 748 169
rect 36 118 41 124
rect 34 117 41 118
rect 34 113 35 117
rect 39 113 41 117
rect 34 112 41 113
rect 43 122 49 124
rect 43 117 51 122
rect 43 113 45 117
rect 49 113 51 117
rect 43 112 51 113
rect 53 117 61 122
rect 53 113 55 117
rect 59 113 61 117
rect 53 112 61 113
rect 63 121 70 122
rect 63 117 65 121
rect 69 117 70 121
rect 122 119 127 140
rect 63 112 70 117
rect 120 118 127 119
rect 120 114 121 118
rect 125 114 127 118
rect 120 113 127 114
rect 129 139 141 140
rect 129 135 131 139
rect 135 135 141 139
rect 129 132 141 135
rect 129 128 131 132
rect 135 131 141 132
rect 158 131 163 140
rect 135 128 143 131
rect 129 113 143 128
rect 145 118 153 131
rect 145 114 147 118
rect 151 114 153 118
rect 145 113 153 114
rect 155 125 163 131
rect 155 121 157 125
rect 161 121 163 125
rect 155 113 163 121
rect 165 134 170 140
rect 165 133 172 134
rect 165 129 167 133
rect 171 129 172 133
rect 165 128 172 129
rect 165 113 170 128
rect 206 119 211 140
rect 204 118 211 119
rect 204 114 205 118
rect 209 114 211 118
rect 204 113 211 114
rect 213 139 225 140
rect 213 135 215 139
rect 219 135 225 139
rect 213 132 225 135
rect 213 128 215 132
rect 219 131 225 132
rect 242 131 247 140
rect 219 128 227 131
rect 213 113 227 128
rect 229 118 237 131
rect 229 114 231 118
rect 235 114 237 118
rect 229 113 237 114
rect 239 125 247 131
rect 239 121 241 125
rect 245 121 247 125
rect 239 113 247 121
rect 249 134 254 140
rect 249 133 256 134
rect 249 129 251 133
rect 255 129 256 133
rect 249 128 256 129
rect 249 113 254 128
rect 268 118 273 124
rect 266 117 273 118
rect 266 113 267 117
rect 271 113 273 117
rect 266 112 273 113
rect 275 122 281 124
rect 275 117 283 122
rect 275 113 277 117
rect 281 113 283 117
rect 275 112 283 113
rect 285 117 293 122
rect 285 113 287 117
rect 291 113 293 117
rect 285 112 293 113
rect 295 121 302 122
rect 295 117 297 121
rect 301 117 302 121
rect 365 120 370 126
rect 295 112 302 117
rect 363 119 370 120
rect 363 115 364 119
rect 368 115 370 119
rect 363 114 370 115
rect 372 124 378 126
rect 372 119 380 124
rect 372 115 374 119
rect 378 115 380 119
rect 372 114 380 115
rect 382 119 390 124
rect 382 115 384 119
rect 388 115 390 119
rect 382 114 390 115
rect 392 123 399 124
rect 392 119 394 123
rect 398 119 399 123
rect 451 121 456 142
rect 392 114 399 119
rect 449 120 456 121
rect 449 116 450 120
rect 454 116 456 120
rect 449 115 456 116
rect 458 141 470 142
rect 458 137 460 141
rect 464 137 470 141
rect 458 134 470 137
rect 458 130 460 134
rect 464 133 470 134
rect 487 133 492 142
rect 464 130 472 133
rect 458 115 472 130
rect 474 120 482 133
rect 474 116 476 120
rect 480 116 482 120
rect 474 115 482 116
rect 484 127 492 133
rect 484 123 486 127
rect 490 123 492 127
rect 484 115 492 123
rect 494 136 499 142
rect 494 135 501 136
rect 494 131 496 135
rect 500 131 501 135
rect 494 130 501 131
rect 494 115 499 130
rect 535 121 540 142
rect 533 120 540 121
rect 533 116 534 120
rect 538 116 540 120
rect 533 115 540 116
rect 542 141 554 142
rect 542 137 544 141
rect 548 137 554 141
rect 542 134 554 137
rect 542 130 544 134
rect 548 133 554 134
rect 571 133 576 142
rect 548 130 556 133
rect 542 115 556 130
rect 558 120 566 133
rect 558 116 560 120
rect 564 116 566 120
rect 558 115 566 116
rect 568 127 576 133
rect 568 123 570 127
rect 574 123 576 127
rect 568 115 576 123
rect 578 136 583 142
rect 578 135 585 136
rect 578 131 580 135
rect 584 131 585 135
rect 578 130 585 131
rect 578 115 583 130
rect 597 120 602 126
rect 595 119 602 120
rect 595 115 596 119
rect 600 115 602 119
rect 595 114 602 115
rect 604 124 610 126
rect 604 119 612 124
rect 604 115 606 119
rect 610 115 612 119
rect 604 114 612 115
rect 614 119 622 124
rect 614 115 616 119
rect 620 115 622 119
rect 614 114 622 115
rect 624 123 631 124
rect 692 123 697 129
rect 624 119 626 123
rect 630 119 631 123
rect 624 114 631 119
rect 690 122 697 123
rect 690 118 691 122
rect 695 118 697 122
rect 690 117 697 118
rect 699 127 705 129
rect 699 122 707 127
rect 699 118 701 122
rect 705 118 707 122
rect 699 117 707 118
rect 709 122 717 127
rect 709 118 711 122
rect 715 118 717 122
rect 709 117 717 118
rect 719 126 726 127
rect 719 122 721 126
rect 725 122 726 126
rect 778 124 783 145
rect 719 117 726 122
rect 776 123 783 124
rect 776 119 777 123
rect 781 119 783 123
rect 776 118 783 119
rect 785 144 797 145
rect 785 140 787 144
rect 791 140 797 144
rect 785 137 797 140
rect 785 133 787 137
rect 791 136 797 137
rect 814 136 819 145
rect 791 133 799 136
rect 785 118 799 133
rect 801 123 809 136
rect 801 119 803 123
rect 807 119 809 123
rect 801 118 809 119
rect 811 130 819 136
rect 811 126 813 130
rect 817 126 819 130
rect 811 118 819 126
rect 821 139 826 145
rect 821 138 828 139
rect 821 134 823 138
rect 827 134 828 138
rect 821 133 828 134
rect 821 118 826 133
rect 862 124 867 145
rect 860 123 867 124
rect 860 119 861 123
rect 865 119 867 123
rect 860 118 867 119
rect 869 144 881 145
rect 869 140 871 144
rect 875 140 881 144
rect 869 137 881 140
rect 869 133 871 137
rect 875 136 881 137
rect 898 136 903 145
rect 875 133 883 136
rect 869 118 883 133
rect 885 123 893 136
rect 885 119 887 123
rect 891 119 893 123
rect 885 118 893 119
rect 895 130 903 136
rect 895 126 897 130
rect 901 126 903 130
rect 895 118 903 126
rect 905 139 910 145
rect 905 138 912 139
rect 905 134 907 138
rect 911 134 912 138
rect 905 133 912 134
rect 905 118 910 133
rect 924 123 929 129
rect 922 122 929 123
rect 922 118 923 122
rect 927 118 929 122
rect 922 117 929 118
rect 931 127 937 129
rect 931 122 939 127
rect 931 118 933 122
rect 937 118 939 122
rect 931 117 939 118
rect 941 122 949 127
rect 941 118 943 122
rect 947 118 949 122
rect 941 117 949 118
rect 951 126 958 127
rect 951 122 953 126
rect 957 122 958 126
rect 951 117 958 122
rect 146 28 154 31
rect 129 23 134 28
rect 127 22 134 23
rect 127 18 128 22
rect 132 18 134 22
rect 127 17 134 18
rect 129 10 134 17
rect 136 10 141 28
rect 143 19 154 28
rect 156 25 161 31
rect 802 33 810 36
rect 475 30 483 33
rect 458 25 463 30
rect 156 24 163 25
rect 156 20 158 24
rect 162 20 163 24
rect 156 19 163 20
rect 456 24 463 25
rect 456 20 457 24
rect 461 20 463 24
rect 456 19 463 20
rect 143 15 152 19
rect 143 11 146 15
rect 150 11 152 15
rect 143 10 152 11
rect 458 12 463 19
rect 465 12 470 30
rect 472 21 483 30
rect 485 27 490 33
rect 785 28 790 33
rect 783 27 790 28
rect 485 26 492 27
rect 485 22 487 26
rect 491 22 492 26
rect 783 23 784 27
rect 788 23 790 27
rect 783 22 790 23
rect 485 21 492 22
rect 472 17 481 21
rect 472 13 475 17
rect 479 13 481 17
rect 785 15 790 22
rect 792 15 797 33
rect 799 24 810 33
rect 812 30 817 36
rect 812 29 819 30
rect 812 25 814 29
rect 818 25 819 29
rect 812 24 819 25
rect 799 20 808 24
rect 799 16 802 20
rect 806 16 808 20
rect 799 15 808 16
rect 472 12 481 13
rect 35 -28 40 -22
rect 33 -29 40 -28
rect 33 -33 34 -29
rect 38 -33 40 -29
rect 33 -34 40 -33
rect 42 -24 48 -22
rect 42 -29 50 -24
rect 42 -33 44 -29
rect 48 -33 50 -29
rect 42 -34 50 -33
rect 52 -29 60 -24
rect 52 -33 54 -29
rect 58 -33 60 -29
rect 52 -34 60 -33
rect 62 -25 69 -24
rect 62 -29 64 -25
rect 68 -29 69 -25
rect 121 -27 126 -6
rect 62 -34 69 -29
rect 119 -28 126 -27
rect 119 -32 120 -28
rect 124 -32 126 -28
rect 119 -33 126 -32
rect 128 -7 140 -6
rect 128 -11 130 -7
rect 134 -11 140 -7
rect 128 -14 140 -11
rect 128 -18 130 -14
rect 134 -15 140 -14
rect 157 -15 162 -6
rect 134 -18 142 -15
rect 128 -33 142 -18
rect 144 -28 152 -15
rect 144 -32 146 -28
rect 150 -32 152 -28
rect 144 -33 152 -32
rect 154 -21 162 -15
rect 154 -25 156 -21
rect 160 -25 162 -21
rect 154 -33 162 -25
rect 164 -12 169 -6
rect 164 -13 171 -12
rect 164 -17 166 -13
rect 170 -17 171 -13
rect 164 -18 171 -17
rect 164 -33 169 -18
rect 205 -27 210 -6
rect 203 -28 210 -27
rect 203 -32 204 -28
rect 208 -32 210 -28
rect 203 -33 210 -32
rect 212 -7 224 -6
rect 212 -11 214 -7
rect 218 -11 224 -7
rect 212 -14 224 -11
rect 212 -18 214 -14
rect 218 -15 224 -14
rect 241 -15 246 -6
rect 218 -18 226 -15
rect 212 -33 226 -18
rect 228 -28 236 -15
rect 228 -32 230 -28
rect 234 -32 236 -28
rect 228 -33 236 -32
rect 238 -21 246 -15
rect 238 -25 240 -21
rect 244 -25 246 -21
rect 238 -33 246 -25
rect 248 -12 253 -6
rect 248 -13 255 -12
rect 248 -17 250 -13
rect 254 -17 255 -13
rect 248 -18 255 -17
rect 248 -33 253 -18
rect 267 -28 272 -22
rect 265 -29 272 -28
rect 265 -33 266 -29
rect 270 -33 272 -29
rect 265 -34 272 -33
rect 274 -24 280 -22
rect 274 -29 282 -24
rect 274 -33 276 -29
rect 280 -33 282 -29
rect 274 -34 282 -33
rect 284 -29 292 -24
rect 284 -33 286 -29
rect 290 -33 292 -29
rect 284 -34 292 -33
rect 294 -25 301 -24
rect 294 -29 296 -25
rect 300 -29 301 -25
rect 364 -26 369 -20
rect 294 -34 301 -29
rect 362 -27 369 -26
rect 362 -31 363 -27
rect 367 -31 369 -27
rect 362 -32 369 -31
rect 371 -22 377 -20
rect 371 -27 379 -22
rect 371 -31 373 -27
rect 377 -31 379 -27
rect 371 -32 379 -31
rect 381 -27 389 -22
rect 381 -31 383 -27
rect 387 -31 389 -27
rect 381 -32 389 -31
rect 391 -23 398 -22
rect 391 -27 393 -23
rect 397 -27 398 -23
rect 450 -25 455 -4
rect 391 -32 398 -27
rect 448 -26 455 -25
rect 448 -30 449 -26
rect 453 -30 455 -26
rect 448 -31 455 -30
rect 457 -5 469 -4
rect 457 -9 459 -5
rect 463 -9 469 -5
rect 457 -12 469 -9
rect 457 -16 459 -12
rect 463 -13 469 -12
rect 486 -13 491 -4
rect 463 -16 471 -13
rect 457 -31 471 -16
rect 473 -26 481 -13
rect 473 -30 475 -26
rect 479 -30 481 -26
rect 473 -31 481 -30
rect 483 -19 491 -13
rect 483 -23 485 -19
rect 489 -23 491 -19
rect 483 -31 491 -23
rect 493 -10 498 -4
rect 493 -11 500 -10
rect 493 -15 495 -11
rect 499 -15 500 -11
rect 493 -16 500 -15
rect 493 -31 498 -16
rect 534 -25 539 -4
rect 532 -26 539 -25
rect 532 -30 533 -26
rect 537 -30 539 -26
rect 532 -31 539 -30
rect 541 -5 553 -4
rect 541 -9 543 -5
rect 547 -9 553 -5
rect 541 -12 553 -9
rect 541 -16 543 -12
rect 547 -13 553 -12
rect 570 -13 575 -4
rect 547 -16 555 -13
rect 541 -31 555 -16
rect 557 -26 565 -13
rect 557 -30 559 -26
rect 563 -30 565 -26
rect 557 -31 565 -30
rect 567 -19 575 -13
rect 567 -23 569 -19
rect 573 -23 575 -19
rect 567 -31 575 -23
rect 577 -10 582 -4
rect 577 -11 584 -10
rect 577 -15 579 -11
rect 583 -15 584 -11
rect 577 -16 584 -15
rect 577 -31 582 -16
rect 596 -26 601 -20
rect 594 -27 601 -26
rect 594 -31 595 -27
rect 599 -31 601 -27
rect 594 -32 601 -31
rect 603 -22 609 -20
rect 603 -27 611 -22
rect 603 -31 605 -27
rect 609 -31 611 -27
rect 603 -32 611 -31
rect 613 -27 621 -22
rect 613 -31 615 -27
rect 619 -31 621 -27
rect 613 -32 621 -31
rect 623 -23 630 -22
rect 691 -23 696 -17
rect 623 -27 625 -23
rect 629 -27 630 -23
rect 623 -32 630 -27
rect 689 -24 696 -23
rect 689 -28 690 -24
rect 694 -28 696 -24
rect 689 -29 696 -28
rect 698 -19 704 -17
rect 698 -24 706 -19
rect 698 -28 700 -24
rect 704 -28 706 -24
rect 698 -29 706 -28
rect 708 -24 716 -19
rect 708 -28 710 -24
rect 714 -28 716 -24
rect 708 -29 716 -28
rect 718 -20 725 -19
rect 718 -24 720 -20
rect 724 -24 725 -20
rect 777 -22 782 -1
rect 718 -29 725 -24
rect 775 -23 782 -22
rect 775 -27 776 -23
rect 780 -27 782 -23
rect 775 -28 782 -27
rect 784 -2 796 -1
rect 784 -6 786 -2
rect 790 -6 796 -2
rect 784 -9 796 -6
rect 784 -13 786 -9
rect 790 -10 796 -9
rect 813 -10 818 -1
rect 790 -13 798 -10
rect 784 -28 798 -13
rect 800 -23 808 -10
rect 800 -27 802 -23
rect 806 -27 808 -23
rect 800 -28 808 -27
rect 810 -16 818 -10
rect 810 -20 812 -16
rect 816 -20 818 -16
rect 810 -28 818 -20
rect 820 -7 825 -1
rect 820 -8 827 -7
rect 820 -12 822 -8
rect 826 -12 827 -8
rect 820 -13 827 -12
rect 820 -28 825 -13
rect 861 -22 866 -1
rect 859 -23 866 -22
rect 859 -27 860 -23
rect 864 -27 866 -23
rect 859 -28 866 -27
rect 868 -2 880 -1
rect 868 -6 870 -2
rect 874 -6 880 -2
rect 868 -9 880 -6
rect 868 -13 870 -9
rect 874 -10 880 -9
rect 897 -10 902 -1
rect 874 -13 882 -10
rect 868 -28 882 -13
rect 884 -23 892 -10
rect 884 -27 886 -23
rect 890 -27 892 -23
rect 884 -28 892 -27
rect 894 -16 902 -10
rect 894 -20 896 -16
rect 900 -20 902 -16
rect 894 -28 902 -20
rect 904 -7 909 -1
rect 904 -8 911 -7
rect 904 -12 906 -8
rect 910 -12 911 -8
rect 904 -13 911 -12
rect 904 -28 909 -13
rect 923 -23 928 -17
rect 921 -24 928 -23
rect 921 -28 922 -24
rect 926 -28 928 -24
rect 921 -29 928 -28
rect 930 -19 936 -17
rect 930 -24 938 -19
rect 930 -28 932 -24
rect 936 -28 938 -24
rect 930 -29 938 -28
rect 940 -24 948 -19
rect 940 -28 942 -24
rect 946 -28 948 -24
rect 940 -29 948 -28
rect 950 -20 957 -19
rect 950 -24 952 -20
rect 956 -24 957 -20
rect 950 -29 957 -24
rect 145 -118 153 -115
rect 128 -123 133 -118
rect 126 -124 133 -123
rect 126 -128 127 -124
rect 131 -128 133 -124
rect 126 -129 133 -128
rect 128 -136 133 -129
rect 135 -136 140 -118
rect 142 -127 153 -118
rect 155 -121 160 -115
rect 801 -113 809 -110
rect 474 -116 482 -113
rect 457 -121 462 -116
rect 155 -122 162 -121
rect 155 -126 157 -122
rect 161 -126 162 -122
rect 155 -127 162 -126
rect 455 -122 462 -121
rect 455 -126 456 -122
rect 460 -126 462 -122
rect 455 -127 462 -126
rect 142 -131 151 -127
rect 142 -135 145 -131
rect 149 -135 151 -131
rect 142 -136 151 -135
rect 457 -134 462 -127
rect 464 -134 469 -116
rect 471 -125 482 -116
rect 484 -119 489 -113
rect 784 -118 789 -113
rect 782 -119 789 -118
rect 484 -120 491 -119
rect 484 -124 486 -120
rect 490 -124 491 -120
rect 782 -123 783 -119
rect 787 -123 789 -119
rect 782 -124 789 -123
rect 484 -125 491 -124
rect 471 -129 480 -125
rect 471 -133 474 -129
rect 478 -133 480 -129
rect 784 -131 789 -124
rect 791 -131 796 -113
rect 798 -122 809 -113
rect 811 -116 816 -110
rect 811 -117 818 -116
rect 811 -121 813 -117
rect 817 -121 818 -117
rect 811 -122 818 -121
rect 798 -126 807 -122
rect 798 -130 801 -126
rect 805 -130 807 -126
rect 798 -131 807 -130
rect 471 -134 480 -133
rect 338 -163 344 -161
rect 329 -168 334 -163
rect 327 -169 334 -168
rect 327 -173 328 -169
rect 332 -173 334 -169
rect 327 -176 334 -173
rect 327 -180 328 -176
rect 332 -180 334 -176
rect 327 -181 334 -180
rect 336 -164 344 -163
rect 336 -168 338 -164
rect 342 -168 344 -164
rect 336 -174 344 -168
rect 346 -162 354 -161
rect 346 -166 348 -162
rect 352 -166 354 -162
rect 346 -169 354 -166
rect 346 -173 348 -169
rect 352 -173 354 -169
rect 346 -174 354 -173
rect 356 -162 363 -161
rect 356 -166 358 -162
rect 362 -166 363 -162
rect 431 -163 437 -161
rect 356 -174 363 -166
rect 422 -168 427 -163
rect 420 -169 427 -168
rect 420 -173 421 -169
rect 425 -173 427 -169
rect 336 -181 342 -174
rect 420 -176 427 -173
rect 420 -180 421 -176
rect 425 -180 427 -176
rect 420 -181 427 -180
rect 429 -164 437 -163
rect 429 -168 431 -164
rect 435 -168 437 -164
rect 429 -174 437 -168
rect 439 -162 447 -161
rect 439 -166 441 -162
rect 445 -166 447 -162
rect 439 -169 447 -166
rect 439 -173 441 -169
rect 445 -173 447 -169
rect 439 -174 447 -173
rect 449 -162 456 -161
rect 449 -166 451 -162
rect 455 -166 456 -162
rect 518 -163 524 -161
rect 449 -174 456 -166
rect 509 -168 514 -163
rect 507 -169 514 -168
rect 507 -173 508 -169
rect 512 -173 514 -169
rect 429 -181 435 -174
rect 507 -176 514 -173
rect 507 -180 508 -176
rect 512 -180 514 -176
rect 507 -181 514 -180
rect 516 -164 524 -163
rect 516 -168 518 -164
rect 522 -168 524 -164
rect 516 -174 524 -168
rect 526 -162 534 -161
rect 526 -166 528 -162
rect 532 -166 534 -162
rect 526 -169 534 -166
rect 526 -173 528 -169
rect 532 -173 534 -169
rect 526 -174 534 -173
rect 536 -162 543 -161
rect 536 -166 538 -162
rect 542 -166 543 -162
rect 536 -174 543 -166
rect 516 -181 522 -174
<< metal1 >>
rect 31 234 472 238
rect 31 212 35 234
rect 113 225 114 228
rect 329 225 522 226
rect 528 225 572 227
rect 113 224 572 225
rect 621 224 665 227
rect 708 226 752 227
rect 708 224 760 226
rect 108 223 760 224
rect 108 221 534 223
rect 108 217 132 221
rect 136 217 142 221
rect 146 217 219 221
rect 223 217 229 221
rect 233 217 312 221
rect 316 217 322 221
rect 326 220 534 221
rect 326 217 332 220
rect 528 219 534 220
rect 538 219 544 223
rect 548 220 627 223
rect 548 219 572 220
rect 621 219 627 220
rect 631 219 637 223
rect 641 220 714 223
rect 641 219 665 220
rect 708 219 714 220
rect 718 219 724 223
rect 728 220 760 223
rect 728 219 752 220
rect 112 207 113 211
rect 117 207 132 211
rect 112 200 124 204
rect 119 195 124 200
rect 128 203 132 207
rect 136 209 148 212
rect 136 206 143 209
rect 147 205 148 209
rect 199 207 200 211
rect 204 207 219 211
rect 143 204 148 205
rect 128 199 140 203
rect 136 195 140 199
rect 119 191 126 195
rect 130 191 133 195
rect 112 178 116 187
rect 120 183 125 187
rect 136 180 140 191
rect 144 190 148 204
rect 200 200 211 204
rect 206 195 211 200
rect 215 203 219 207
rect 223 209 235 212
rect 223 206 230 209
rect 234 205 235 209
rect 292 207 293 211
rect 297 207 312 211
rect 230 204 235 205
rect 215 199 227 203
rect 223 195 227 199
rect 206 191 213 195
rect 217 191 220 195
rect 144 187 173 190
rect 144 186 148 187
rect 105 174 116 178
rect 123 178 140 180
rect 127 176 140 178
rect 143 185 148 186
rect 147 181 148 185
rect 143 178 148 181
rect 123 171 127 174
rect 147 174 148 178
rect 143 173 148 174
rect 112 167 113 171
rect 117 167 118 171
rect 112 161 118 167
rect 123 166 127 167
rect 132 169 133 173
rect 137 169 138 173
rect 132 161 138 169
rect 108 157 142 161
rect 146 157 152 161
rect 108 153 152 157
rect 109 146 113 153
rect 169 151 173 187
rect 199 177 203 187
rect 207 183 212 187
rect 223 180 227 191
rect 231 186 235 204
rect 293 200 304 204
rect 299 195 304 200
rect 308 203 312 207
rect 316 209 328 212
rect 532 211 544 214
rect 316 206 323 209
rect 327 205 328 209
rect 341 205 513 209
rect 518 205 519 209
rect 532 207 533 211
rect 537 208 544 211
rect 548 209 563 213
rect 567 209 568 213
rect 625 211 637 214
rect 532 206 537 207
rect 323 204 328 205
rect 308 199 320 203
rect 316 195 320 199
rect 299 191 306 195
rect 310 191 313 195
rect 196 174 203 177
rect 210 178 227 180
rect 214 176 227 178
rect 230 185 235 186
rect 234 181 235 185
rect 230 178 235 181
rect 210 171 214 174
rect 234 176 235 178
rect 234 174 241 176
rect 230 173 241 174
rect 292 177 296 187
rect 300 183 305 187
rect 316 180 320 191
rect 324 186 328 204
rect 532 199 536 206
rect 548 205 552 209
rect 625 207 626 211
rect 630 208 637 211
rect 641 209 656 213
rect 660 209 661 213
rect 712 211 724 214
rect 625 206 630 207
rect 476 195 536 199
rect 532 188 536 195
rect 540 201 552 205
rect 556 203 567 206
rect 540 197 544 201
rect 556 197 561 203
rect 547 193 550 197
rect 554 193 561 197
rect 625 195 629 206
rect 641 205 645 209
rect 712 207 713 211
rect 717 208 724 211
rect 728 209 743 213
rect 747 209 748 213
rect 712 206 717 207
rect 532 187 537 188
rect 289 174 296 177
rect 303 178 320 180
rect 307 176 320 178
rect 323 185 328 186
rect 327 181 328 185
rect 341 183 514 186
rect 532 183 533 187
rect 323 178 328 181
rect 199 167 200 171
rect 204 167 205 171
rect 199 161 205 167
rect 210 166 214 167
rect 219 169 220 173
rect 224 169 225 173
rect 303 171 307 174
rect 327 174 328 178
rect 532 180 537 183
rect 532 176 533 180
rect 540 182 544 193
rect 602 192 629 195
rect 555 185 560 189
rect 540 180 557 182
rect 540 178 553 180
rect 532 175 537 176
rect 564 179 568 189
rect 602 180 606 192
rect 564 176 571 179
rect 323 173 328 174
rect 219 161 225 169
rect 292 167 293 171
rect 297 167 298 171
rect 292 161 298 167
rect 303 166 307 167
rect 312 169 313 173
rect 317 169 318 173
rect 542 171 543 175
rect 547 171 548 175
rect 312 161 318 169
rect 341 165 515 168
rect 542 163 548 171
rect 553 173 557 176
rect 625 188 629 192
rect 633 201 645 205
rect 649 205 663 206
rect 649 203 660 205
rect 633 197 637 201
rect 649 197 654 203
rect 640 193 643 197
rect 647 193 654 197
rect 625 187 630 188
rect 625 183 626 187
rect 625 180 630 183
rect 625 176 626 180
rect 633 182 637 193
rect 712 192 716 206
rect 728 205 732 209
rect 648 185 653 189
rect 633 180 650 182
rect 633 178 646 180
rect 625 175 630 176
rect 657 179 661 189
rect 690 188 716 192
rect 720 201 732 205
rect 736 205 750 206
rect 736 203 747 205
rect 720 197 724 201
rect 736 197 741 203
rect 727 193 730 197
rect 734 193 741 197
rect 657 176 664 179
rect 676 178 677 182
rect 553 168 557 169
rect 562 169 563 173
rect 567 169 568 173
rect 562 163 568 169
rect 635 171 636 175
rect 640 171 641 175
rect 635 163 641 171
rect 646 173 650 176
rect 646 168 650 169
rect 655 169 656 173
rect 660 169 661 173
rect 655 163 661 169
rect 195 157 229 161
rect 233 157 239 161
rect 195 156 239 157
rect 288 157 322 161
rect 326 157 332 161
rect 195 153 222 156
rect 288 153 332 157
rect 528 159 534 163
rect 538 159 572 163
rect 621 159 627 163
rect 631 159 665 163
rect 528 155 572 159
rect 197 146 201 153
rect 234 149 267 152
rect 288 146 292 153
rect 564 151 568 155
rect 583 154 613 157
rect 621 155 665 159
rect 676 158 680 178
rect 522 150 626 151
rect 522 148 648 150
rect 657 148 661 155
rect 690 157 694 188
rect 712 187 717 188
rect 712 183 713 187
rect 700 158 704 178
rect 712 180 717 183
rect 712 176 713 180
rect 720 182 724 193
rect 735 185 740 189
rect 720 180 737 182
rect 720 178 733 180
rect 712 175 717 176
rect 744 180 748 189
rect 744 176 752 180
rect 722 171 723 175
rect 727 171 728 175
rect 722 163 728 171
rect 733 173 737 176
rect 733 168 737 169
rect 742 169 743 173
rect 747 169 748 173
rect 742 163 748 169
rect 708 159 714 163
rect 718 159 752 163
rect 708 155 752 159
rect 746 148 750 155
rect 760 148 962 151
rect 304 147 962 148
rect 304 146 692 147
rect 0 145 227 146
rect 240 145 692 146
rect 0 144 692 145
rect 0 142 365 144
rect 0 138 36 142
rect 40 138 50 142
rect 54 138 64 142
rect 68 139 147 142
rect 68 138 131 139
rect 0 27 4 138
rect 20 137 35 138
rect 34 118 38 125
rect 34 117 39 118
rect 34 113 35 117
rect 42 117 46 138
rect 49 132 62 133
rect 49 128 52 132
rect 56 128 58 132
rect 49 127 62 128
rect 49 120 55 127
rect 65 121 69 138
rect 135 138 147 139
rect 151 139 231 142
rect 151 138 215 139
rect 112 127 124 133
rect 131 132 135 135
rect 219 138 231 139
rect 235 138 268 142
rect 272 138 282 142
rect 286 138 296 142
rect 300 140 365 142
rect 369 140 379 144
rect 383 140 393 144
rect 397 141 476 144
rect 397 140 460 141
rect 300 138 335 140
rect 145 129 167 133
rect 171 129 172 133
rect 196 132 208 133
rect 145 128 149 129
rect 131 127 135 128
rect 112 124 117 127
rect 112 123 113 124
rect 42 113 45 117
rect 49 113 50 117
rect 54 113 55 117
rect 59 113 60 117
rect 65 116 69 117
rect 104 120 113 123
rect 138 124 149 128
rect 196 128 201 132
rect 205 128 208 132
rect 196 127 208 128
rect 215 132 219 135
rect 229 129 251 133
rect 255 129 256 133
rect 229 128 233 129
rect 215 127 219 128
rect 138 120 142 124
rect 156 121 157 125
rect 161 121 172 125
rect 34 112 39 113
rect 34 104 38 112
rect 54 108 60 113
rect 41 104 42 108
rect 46 104 60 108
rect 66 106 70 109
rect 104 106 107 120
rect 112 119 117 120
rect 121 118 142 120
rect 34 95 38 100
rect 34 94 39 95
rect 34 90 35 94
rect 39 90 46 93
rect 34 87 46 90
rect 50 91 54 104
rect 113 114 121 115
rect 125 116 142 118
rect 113 111 125 114
rect 66 100 70 102
rect 57 96 61 100
rect 65 96 70 100
rect 57 95 70 96
rect 113 99 117 111
rect 138 109 142 116
rect 146 114 147 118
rect 151 117 152 118
rect 151 114 163 117
rect 146 113 163 114
rect 159 110 163 113
rect 159 109 164 110
rect 127 103 133 108
rect 138 105 150 109
rect 154 105 155 109
rect 159 105 160 109
rect 127 101 129 103
rect 120 99 129 101
rect 159 104 164 105
rect 168 105 172 121
rect 196 124 201 127
rect 196 120 197 124
rect 222 124 233 128
rect 222 120 226 124
rect 240 121 241 125
rect 245 121 256 125
rect 196 119 201 120
rect 205 118 226 120
rect 197 114 205 115
rect 209 116 226 118
rect 197 111 209 114
rect 159 100 163 104
rect 120 95 133 99
rect 139 96 163 100
rect 168 101 170 105
rect 113 94 117 95
rect 139 94 143 96
rect 50 87 64 91
rect 68 87 69 91
rect 126 87 127 91
rect 131 87 132 91
rect 168 92 172 101
rect 197 99 201 111
rect 222 109 226 116
rect 230 114 231 118
rect 235 117 236 118
rect 235 114 247 117
rect 230 113 247 114
rect 243 110 247 113
rect 243 109 248 110
rect 211 103 217 108
rect 222 105 234 109
rect 238 105 239 109
rect 243 105 244 109
rect 211 101 213 103
rect 204 99 213 101
rect 243 104 248 105
rect 243 100 247 104
rect 204 95 217 99
rect 223 96 247 100
rect 197 94 201 95
rect 223 94 227 96
rect 139 89 143 90
rect 148 88 149 92
rect 153 88 172 92
rect 126 82 132 87
rect 210 87 211 91
rect 215 87 216 91
rect 252 92 256 121
rect 266 118 270 125
rect 266 117 271 118
rect 266 113 267 117
rect 274 117 278 138
rect 281 132 294 133
rect 281 128 284 132
rect 288 128 290 132
rect 281 127 294 128
rect 281 120 287 127
rect 297 121 301 138
rect 274 113 277 117
rect 281 113 282 117
rect 286 113 287 117
rect 291 113 292 117
rect 297 116 301 117
rect 266 112 271 113
rect 266 104 270 112
rect 286 108 292 113
rect 273 104 274 108
rect 278 104 292 108
rect 298 107 302 109
rect 223 89 227 90
rect 232 88 233 92
rect 237 88 256 92
rect 260 101 270 104
rect 260 89 263 101
rect 210 82 216 87
rect 266 95 270 101
rect 266 94 271 95
rect 266 90 267 94
rect 271 90 278 93
rect 266 87 278 90
rect 282 91 286 104
rect 298 100 302 103
rect 289 96 293 100
rect 297 96 302 100
rect 289 95 302 96
rect 282 87 296 91
rect 300 87 301 91
rect 33 78 36 82
rect 40 78 46 82
rect 50 78 114 82
rect 118 78 167 82
rect 171 78 198 82
rect 202 78 251 82
rect 255 78 268 82
rect 272 78 278 82
rect 282 81 306 82
rect 282 78 300 81
rect 19 75 300 78
rect 19 74 306 75
rect 123 72 167 74
rect 123 68 129 72
rect 133 68 157 72
rect 161 68 167 72
rect 127 60 133 68
rect 127 56 128 60
rect 132 56 133 60
rect 138 60 142 61
rect 147 60 153 68
rect 147 56 148 60
rect 152 56 153 60
rect 158 60 163 63
rect 162 56 163 60
rect 138 53 142 56
rect 158 55 163 56
rect 138 49 155 53
rect 127 37 131 47
rect 135 42 140 46
rect 151 45 155 49
rect 135 34 141 38
rect 145 34 148 38
rect -1 7 4 27
rect 135 28 139 34
rect 151 30 155 41
rect 122 25 139 28
rect 143 26 155 30
rect 159 51 320 55
rect 143 22 147 26
rect 159 25 163 51
rect 329 29 333 138
rect 363 120 367 127
rect 363 119 368 120
rect 363 115 364 119
rect 371 119 375 140
rect 378 134 391 135
rect 378 130 381 134
rect 385 130 387 134
rect 378 129 391 130
rect 378 122 384 129
rect 394 123 398 140
rect 464 140 476 141
rect 480 141 560 144
rect 480 140 544 141
rect 441 129 453 135
rect 460 134 464 137
rect 548 140 560 141
rect 564 140 597 144
rect 601 140 611 144
rect 615 140 625 144
rect 629 143 692 144
rect 696 143 706 147
rect 710 143 720 147
rect 724 144 803 147
rect 724 143 787 144
rect 629 140 665 143
rect 474 131 496 135
rect 500 131 501 135
rect 516 134 537 135
rect 474 130 478 131
rect 460 129 464 130
rect 441 126 446 129
rect 441 125 442 126
rect 371 115 374 119
rect 378 115 379 119
rect 383 115 384 119
rect 388 115 389 119
rect 394 118 398 119
rect 433 122 442 125
rect 467 126 478 130
rect 516 130 530 134
rect 534 130 537 134
rect 516 129 537 130
rect 544 134 548 137
rect 558 131 580 135
rect 584 131 585 135
rect 558 130 562 131
rect 544 129 548 130
rect 467 122 471 126
rect 485 123 486 127
rect 490 123 501 127
rect 363 114 368 115
rect 363 106 367 114
rect 383 110 389 115
rect 370 106 371 110
rect 375 106 389 110
rect 395 108 399 111
rect 433 108 436 122
rect 441 121 446 122
rect 450 120 471 122
rect 363 97 367 102
rect 363 96 368 97
rect 363 92 364 96
rect 368 92 375 95
rect 363 89 375 92
rect 379 93 383 106
rect 442 116 450 117
rect 454 118 471 120
rect 442 113 454 116
rect 395 102 399 104
rect 386 98 390 102
rect 394 98 399 102
rect 386 97 399 98
rect 442 101 446 113
rect 467 111 471 118
rect 475 116 476 120
rect 480 119 481 120
rect 480 116 492 119
rect 475 115 492 116
rect 488 112 492 115
rect 488 111 493 112
rect 456 105 462 110
rect 467 107 479 111
rect 483 107 484 111
rect 488 107 489 111
rect 456 103 458 105
rect 449 101 458 103
rect 488 106 493 107
rect 497 107 501 123
rect 525 126 530 129
rect 525 122 526 126
rect 551 126 562 130
rect 551 122 555 126
rect 569 123 570 127
rect 574 123 587 127
rect 525 121 530 122
rect 534 120 555 122
rect 526 116 534 117
rect 538 118 555 120
rect 526 113 538 116
rect 488 102 492 106
rect 449 97 462 101
rect 468 98 492 102
rect 497 103 499 107
rect 442 96 446 97
rect 468 96 472 98
rect 379 89 393 93
rect 397 89 398 93
rect 455 89 456 93
rect 460 89 461 93
rect 497 94 501 103
rect 526 101 530 113
rect 551 111 555 118
rect 559 116 560 120
rect 564 119 565 120
rect 564 116 576 119
rect 559 115 576 116
rect 572 112 576 115
rect 572 111 577 112
rect 540 105 546 110
rect 551 107 563 111
rect 567 107 568 111
rect 572 107 573 111
rect 540 103 542 105
rect 533 101 542 103
rect 572 106 577 107
rect 572 102 576 106
rect 533 97 546 101
rect 552 98 576 102
rect 526 96 530 97
rect 552 96 556 98
rect 468 91 472 92
rect 477 90 478 94
rect 482 90 501 94
rect 455 84 461 89
rect 539 89 540 93
rect 544 89 545 93
rect 581 94 585 123
rect 595 120 599 127
rect 595 119 600 120
rect 595 115 596 119
rect 603 119 607 140
rect 610 134 623 135
rect 610 130 613 134
rect 617 130 619 134
rect 610 129 623 130
rect 610 122 616 129
rect 626 123 630 140
rect 603 115 606 119
rect 610 115 611 119
rect 615 115 616 119
rect 620 115 621 119
rect 626 118 630 119
rect 595 114 600 115
rect 595 106 599 114
rect 615 110 621 115
rect 602 106 603 110
rect 607 106 621 110
rect 627 109 631 111
rect 552 91 556 92
rect 561 90 562 94
rect 566 90 585 94
rect 589 103 599 106
rect 589 91 592 103
rect 539 84 545 89
rect 595 97 599 103
rect 595 96 600 97
rect 595 92 596 96
rect 600 92 607 95
rect 595 89 607 92
rect 611 93 615 106
rect 627 102 631 105
rect 618 98 622 102
rect 626 98 631 102
rect 618 97 631 98
rect 611 89 625 93
rect 629 89 630 93
rect 362 80 365 84
rect 369 80 375 84
rect 379 80 443 84
rect 447 80 496 84
rect 500 80 527 84
rect 531 80 580 84
rect 584 80 597 84
rect 601 80 607 84
rect 611 83 635 84
rect 611 80 627 83
rect 362 79 627 80
rect 347 77 627 79
rect 633 77 635 83
rect 347 76 635 77
rect 347 75 363 76
rect 452 74 496 76
rect 452 70 458 74
rect 462 70 486 74
rect 490 70 496 74
rect 456 62 462 70
rect 456 58 457 62
rect 461 58 462 62
rect 467 62 471 63
rect 476 62 482 70
rect 476 58 477 62
rect 481 58 482 62
rect 487 62 492 65
rect 491 58 492 62
rect 467 55 471 58
rect 487 57 492 58
rect 349 51 417 55
rect 467 51 484 55
rect 456 39 460 49
rect 464 44 469 48
rect 480 47 484 51
rect 464 36 470 40
rect 474 36 477 40
rect 158 24 163 25
rect 127 18 128 22
rect 132 18 147 22
rect 150 20 158 22
rect 162 20 163 24
rect 150 18 163 20
rect 145 12 146 15
rect 123 11 146 12
rect 150 12 151 15
rect 150 11 157 12
rect 123 8 157 11
rect 161 8 167 12
rect 123 7 167 8
rect 328 9 333 29
rect 464 30 468 36
rect 480 32 484 43
rect 451 27 468 30
rect 472 28 484 32
rect 488 51 492 57
rect 488 48 639 51
rect 643 48 644 51
rect 472 24 476 28
rect 488 27 492 48
rect 656 32 660 140
rect 690 123 694 130
rect 690 122 695 123
rect 690 118 691 122
rect 698 122 702 143
rect 705 137 718 138
rect 705 133 708 137
rect 712 133 714 137
rect 705 132 718 133
rect 705 125 711 132
rect 721 126 725 143
rect 791 143 803 144
rect 807 144 887 147
rect 807 143 871 144
rect 768 132 780 138
rect 787 137 791 140
rect 875 143 887 144
rect 891 143 924 147
rect 928 143 938 147
rect 942 143 952 147
rect 956 143 962 147
rect 801 134 823 138
rect 827 134 828 138
rect 841 137 864 138
rect 801 133 805 134
rect 841 133 857 137
rect 861 133 864 137
rect 787 132 791 133
rect 768 129 773 132
rect 768 128 769 129
rect 698 118 701 122
rect 705 118 706 122
rect 710 118 711 122
rect 715 118 716 122
rect 721 121 725 122
rect 690 117 695 118
rect 690 109 694 117
rect 710 113 716 118
rect 697 109 698 113
rect 702 109 716 113
rect 722 111 726 114
rect 690 100 694 105
rect 690 99 695 100
rect 690 95 691 99
rect 695 95 702 98
rect 690 92 702 95
rect 706 96 710 109
rect 722 105 726 107
rect 713 101 717 105
rect 721 101 726 105
rect 713 100 726 101
rect 706 92 720 96
rect 724 92 725 96
rect 749 94 753 123
rect 760 125 769 128
rect 794 129 805 133
rect 794 125 798 129
rect 812 126 813 130
rect 817 126 828 130
rect 760 111 763 125
rect 768 124 773 125
rect 777 123 798 125
rect 769 119 777 120
rect 781 121 798 123
rect 769 116 781 119
rect 769 104 773 116
rect 794 114 798 121
rect 802 119 803 123
rect 807 122 808 123
rect 807 119 819 122
rect 802 118 819 119
rect 815 115 819 118
rect 815 114 820 115
rect 783 108 789 113
rect 794 110 806 114
rect 810 110 811 114
rect 815 110 816 114
rect 783 106 785 108
rect 776 104 785 106
rect 815 109 820 110
rect 824 110 828 126
rect 815 105 819 109
rect 776 100 789 104
rect 795 101 819 105
rect 824 106 826 110
rect 769 99 773 100
rect 795 99 799 101
rect 749 90 750 94
rect 782 92 783 96
rect 787 92 788 96
rect 824 97 828 106
rect 795 94 799 95
rect 804 93 805 97
rect 809 93 828 97
rect 835 94 838 125
rect 782 87 788 92
rect 842 87 846 133
rect 852 132 864 133
rect 871 137 875 140
rect 885 134 907 138
rect 911 134 912 138
rect 885 133 889 134
rect 871 132 875 133
rect 852 129 857 132
rect 852 125 853 129
rect 878 129 889 133
rect 878 125 882 129
rect 896 126 897 130
rect 901 126 912 130
rect 852 124 857 125
rect 861 123 882 125
rect 853 119 861 120
rect 865 121 882 123
rect 853 116 865 119
rect 853 104 857 116
rect 878 114 882 121
rect 886 119 887 123
rect 891 122 892 123
rect 891 119 903 122
rect 886 118 903 119
rect 899 115 903 118
rect 899 114 904 115
rect 867 108 873 113
rect 878 110 890 114
rect 894 110 895 114
rect 899 110 900 114
rect 867 106 869 108
rect 860 104 869 106
rect 899 109 904 110
rect 899 105 903 109
rect 860 100 873 104
rect 879 101 903 105
rect 853 99 857 100
rect 879 99 883 101
rect 866 92 867 96
rect 871 92 872 96
rect 908 97 912 126
rect 922 123 926 130
rect 922 122 927 123
rect 922 118 923 122
rect 930 122 934 143
rect 937 137 950 138
rect 937 133 940 137
rect 944 133 946 137
rect 937 132 950 133
rect 937 125 943 132
rect 953 126 957 143
rect 930 118 933 122
rect 937 118 938 122
rect 942 118 943 122
rect 947 118 948 122
rect 953 121 957 122
rect 922 117 927 118
rect 922 109 926 117
rect 942 113 948 118
rect 929 109 930 113
rect 934 109 948 113
rect 954 112 958 114
rect 879 94 883 95
rect 888 93 889 97
rect 893 93 912 97
rect 916 106 926 109
rect 916 94 919 106
rect 866 87 872 92
rect 922 100 926 106
rect 922 99 927 100
rect 922 95 923 99
rect 927 95 934 98
rect 922 92 934 95
rect 938 96 942 109
rect 954 105 958 108
rect 945 101 949 105
rect 953 101 958 105
rect 945 100 958 101
rect 938 92 952 96
rect 956 92 957 96
rect 689 86 692 87
rect 687 83 692 86
rect 696 83 702 87
rect 706 83 770 87
rect 774 83 823 87
rect 827 83 854 87
rect 858 83 907 87
rect 911 83 924 87
rect 928 83 934 87
rect 938 83 962 87
rect 687 81 962 83
rect 674 79 962 81
rect 674 78 691 79
rect 674 77 690 78
rect 779 77 823 79
rect 779 73 785 77
rect 789 73 813 77
rect 817 73 823 77
rect 783 65 789 73
rect 783 61 784 65
rect 788 61 789 65
rect 794 65 798 66
rect 803 65 809 73
rect 803 61 804 65
rect 808 61 809 65
rect 814 65 819 68
rect 818 61 819 65
rect 675 48 742 51
rect 746 48 747 51
rect 487 26 492 27
rect 456 20 457 24
rect 461 20 476 24
rect 479 22 487 24
rect 491 22 492 26
rect 479 20 492 22
rect 474 14 475 17
rect 452 13 475 14
rect 479 14 480 17
rect 479 13 486 14
rect 452 10 486 13
rect 490 10 496 14
rect 452 9 496 10
rect -1 4 167 7
rect -1 3 127 4
rect 305 3 320 7
rect 124 0 127 3
rect 328 6 496 9
rect 655 12 660 32
rect 752 20 756 60
rect 794 58 798 61
rect 814 60 819 61
rect 794 54 811 58
rect 764 26 767 53
rect 783 42 787 52
rect 791 47 796 51
rect 807 50 811 54
rect 791 39 797 43
rect 801 39 804 43
rect 791 33 795 39
rect 807 35 811 46
rect 778 30 795 33
rect 799 31 811 35
rect 815 56 819 60
rect 815 53 827 56
rect 799 27 803 31
rect 815 30 819 53
rect 835 32 838 47
rect 814 29 819 30
rect 783 23 784 27
rect 788 23 803 27
rect 806 25 814 27
rect 818 25 819 29
rect 806 23 819 25
rect 801 17 802 20
rect 752 15 756 16
rect 779 16 802 17
rect 806 17 807 20
rect 834 19 839 32
rect 806 16 813 17
rect 779 13 813 16
rect 817 13 823 17
rect 779 12 823 13
rect 655 9 823 12
rect 655 8 779 9
rect 328 5 454 6
rect 784 5 787 9
rect 451 2 454 5
rect -1 -4 305 0
rect -1 -8 35 -4
rect 39 -8 49 -4
rect 53 -8 63 -4
rect 67 -7 146 -4
rect 67 -8 130 -7
rect -1 -119 3 -8
rect 33 -28 37 -21
rect 33 -29 38 -28
rect 33 -33 34 -29
rect 41 -29 45 -8
rect 48 -14 61 -13
rect 48 -18 51 -14
rect 55 -18 57 -14
rect 48 -19 61 -18
rect 48 -26 54 -19
rect 64 -25 68 -8
rect 134 -8 146 -7
rect 150 -7 230 -4
rect 150 -8 214 -7
rect 111 -19 123 -13
rect 130 -14 134 -11
rect 218 -8 230 -7
rect 234 -8 267 -4
rect 271 -8 281 -4
rect 285 -8 295 -4
rect 299 -8 305 -4
rect 328 -2 634 2
rect 328 -6 364 -2
rect 368 -6 378 -2
rect 382 -6 392 -2
rect 396 -5 475 -2
rect 396 -6 459 -5
rect 144 -17 166 -13
rect 170 -17 171 -13
rect 195 -14 207 -13
rect 183 -17 200 -14
rect 144 -18 148 -17
rect 130 -19 134 -18
rect 111 -22 116 -19
rect 111 -23 112 -22
rect 41 -33 44 -29
rect 48 -33 49 -29
rect 53 -33 54 -29
rect 58 -33 59 -29
rect 64 -30 68 -29
rect 103 -26 112 -23
rect 137 -22 148 -18
rect 137 -26 141 -22
rect 155 -25 156 -21
rect 160 -25 171 -21
rect 33 -34 38 -33
rect 33 -42 37 -34
rect 53 -38 59 -33
rect 40 -42 41 -38
rect 45 -42 59 -38
rect 65 -40 69 -37
rect 103 -40 106 -26
rect 111 -27 116 -26
rect 120 -28 141 -26
rect 33 -51 37 -46
rect 33 -52 38 -51
rect 33 -56 34 -52
rect 38 -56 45 -53
rect 33 -59 45 -56
rect 49 -55 53 -42
rect 112 -32 120 -31
rect 124 -30 141 -28
rect 112 -35 124 -32
rect 65 -46 69 -44
rect 56 -50 60 -46
rect 64 -50 69 -46
rect 56 -51 69 -50
rect 112 -47 116 -35
rect 137 -37 141 -30
rect 145 -32 146 -28
rect 150 -29 151 -28
rect 150 -32 162 -29
rect 145 -33 162 -32
rect 158 -36 162 -33
rect 158 -37 163 -36
rect 126 -43 132 -38
rect 137 -41 149 -37
rect 153 -41 154 -37
rect 158 -41 159 -37
rect 126 -45 128 -43
rect 119 -47 128 -45
rect 158 -42 163 -41
rect 167 -41 171 -25
rect 158 -46 162 -42
rect 119 -51 132 -47
rect 138 -50 162 -46
rect 167 -45 169 -41
rect 112 -52 116 -51
rect 138 -52 142 -50
rect 49 -59 63 -55
rect 67 -59 68 -55
rect 125 -59 126 -55
rect 130 -59 131 -55
rect 167 -54 171 -45
rect 138 -57 142 -56
rect 147 -58 148 -54
rect 152 -58 171 -54
rect 183 -57 186 -17
rect 195 -18 200 -17
rect 204 -18 207 -14
rect 195 -19 207 -18
rect 214 -14 218 -11
rect 228 -17 250 -13
rect 254 -17 255 -13
rect 228 -18 232 -17
rect 214 -19 218 -18
rect 195 -22 200 -19
rect 195 -26 196 -22
rect 221 -22 232 -18
rect 221 -26 225 -22
rect 239 -25 240 -21
rect 244 -25 255 -21
rect 195 -27 200 -26
rect 204 -28 225 -26
rect 196 -32 204 -31
rect 208 -30 225 -28
rect 196 -35 208 -32
rect 196 -47 200 -35
rect 221 -37 225 -30
rect 229 -32 230 -28
rect 234 -29 235 -28
rect 234 -32 246 -29
rect 229 -33 246 -32
rect 242 -36 246 -33
rect 242 -37 247 -36
rect 210 -43 216 -38
rect 221 -41 233 -37
rect 237 -41 238 -37
rect 242 -41 243 -37
rect 210 -45 212 -43
rect 203 -47 212 -45
rect 242 -42 247 -41
rect 242 -46 246 -42
rect 203 -51 216 -47
rect 222 -50 246 -46
rect 196 -52 200 -51
rect 222 -52 226 -50
rect 125 -64 131 -59
rect 209 -59 210 -55
rect 214 -59 215 -55
rect 251 -54 255 -25
rect 265 -28 269 -21
rect 265 -29 270 -28
rect 265 -33 266 -29
rect 273 -29 277 -8
rect 280 -14 293 -13
rect 280 -18 283 -14
rect 287 -18 289 -14
rect 280 -19 293 -18
rect 280 -26 286 -19
rect 296 -25 300 -8
rect 273 -33 276 -29
rect 280 -33 281 -29
rect 285 -33 286 -29
rect 290 -33 291 -29
rect 296 -30 300 -29
rect 265 -34 270 -33
rect 265 -42 269 -34
rect 285 -38 291 -33
rect 272 -42 273 -38
rect 277 -42 291 -38
rect 297 -39 301 -37
rect 222 -57 226 -56
rect 231 -58 232 -54
rect 236 -58 255 -54
rect 259 -45 269 -42
rect 259 -57 262 -45
rect 209 -64 215 -59
rect 265 -51 269 -45
rect 265 -52 270 -51
rect 265 -56 266 -52
rect 270 -56 277 -53
rect 265 -59 277 -56
rect 281 -55 285 -42
rect 297 -46 301 -43
rect 288 -50 292 -46
rect 296 -50 301 -46
rect 288 -51 301 -50
rect 281 -59 295 -55
rect 299 -59 300 -55
rect 32 -68 35 -64
rect 39 -68 45 -64
rect 49 -68 113 -64
rect 117 -68 166 -64
rect 170 -68 197 -64
rect 201 -68 250 -64
rect 254 -68 267 -64
rect 271 -68 277 -64
rect 281 -68 300 -64
rect 32 -71 300 -68
rect 32 -72 305 -71
rect 122 -74 166 -72
rect 122 -78 128 -74
rect 132 -78 156 -74
rect 160 -78 166 -74
rect 126 -86 132 -78
rect 126 -90 127 -86
rect 131 -90 132 -86
rect 137 -86 141 -85
rect 146 -86 152 -78
rect 253 -81 294 -78
rect 146 -90 147 -86
rect 151 -90 152 -86
rect 157 -86 162 -83
rect 161 -90 162 -86
rect 137 -93 141 -90
rect 157 -91 162 -90
rect 137 -97 154 -93
rect 126 -109 130 -99
rect 134 -104 139 -100
rect 150 -101 154 -97
rect 134 -112 140 -108
rect 144 -112 147 -108
rect -2 -139 3 -119
rect 134 -118 138 -112
rect 150 -116 154 -105
rect 121 -121 138 -118
rect 142 -120 154 -116
rect 142 -124 146 -120
rect 158 -121 162 -91
rect 250 -99 273 -96
rect 278 -99 279 -96
rect 157 -122 162 -121
rect 126 -128 127 -124
rect 131 -128 146 -124
rect 149 -126 157 -124
rect 161 -126 162 -122
rect 149 -128 162 -126
rect 144 -134 145 -131
rect 122 -135 145 -134
rect 149 -134 150 -131
rect 149 -135 156 -134
rect 122 -138 156 -135
rect 160 -138 166 -134
rect 122 -139 166 -138
rect -2 -142 166 -139
rect -2 -143 122 -142
rect 291 -182 294 -81
rect 303 -100 319 -96
rect 328 -117 332 -6
rect 362 -26 366 -19
rect 362 -27 367 -26
rect 362 -31 363 -27
rect 370 -27 374 -6
rect 377 -12 390 -11
rect 377 -16 380 -12
rect 384 -16 386 -12
rect 377 -17 390 -16
rect 377 -24 383 -17
rect 393 -23 397 -6
rect 463 -6 475 -5
rect 479 -5 559 -2
rect 479 -6 543 -5
rect 440 -17 452 -11
rect 459 -12 463 -9
rect 547 -6 559 -5
rect 563 -6 596 -2
rect 600 -6 610 -2
rect 614 -6 624 -2
rect 628 -6 634 -2
rect 655 1 961 5
rect 655 -3 691 1
rect 695 -3 705 1
rect 709 -3 719 1
rect 723 -2 802 1
rect 723 -3 786 -2
rect 473 -15 495 -11
rect 499 -15 500 -11
rect 524 -12 536 -11
rect 473 -16 477 -15
rect 459 -17 463 -16
rect 440 -20 445 -17
rect 440 -21 441 -20
rect 370 -31 373 -27
rect 377 -31 378 -27
rect 382 -31 383 -27
rect 387 -31 388 -27
rect 393 -28 397 -27
rect 432 -24 441 -21
rect 466 -20 477 -16
rect 524 -16 529 -12
rect 533 -16 536 -12
rect 524 -17 536 -16
rect 543 -12 547 -9
rect 557 -15 579 -11
rect 583 -15 584 -11
rect 557 -16 561 -15
rect 543 -17 547 -16
rect 466 -24 470 -20
rect 484 -23 485 -19
rect 489 -23 500 -19
rect 362 -32 367 -31
rect 362 -40 366 -32
rect 382 -36 388 -31
rect 369 -40 370 -36
rect 374 -40 388 -36
rect 394 -38 398 -35
rect 362 -49 366 -44
rect 362 -50 367 -49
rect 362 -54 363 -50
rect 367 -54 374 -51
rect 362 -57 374 -54
rect 378 -53 382 -40
rect 394 -44 398 -42
rect 385 -48 389 -44
rect 393 -48 398 -44
rect 385 -49 398 -48
rect 378 -57 392 -53
rect 396 -57 397 -53
rect 422 -55 425 -35
rect 432 -38 435 -24
rect 440 -25 445 -24
rect 449 -26 470 -24
rect 441 -30 449 -29
rect 453 -28 470 -26
rect 441 -33 453 -30
rect 441 -45 445 -33
rect 466 -35 470 -28
rect 474 -30 475 -26
rect 479 -27 480 -26
rect 479 -30 491 -27
rect 474 -31 491 -30
rect 487 -34 491 -31
rect 487 -35 492 -34
rect 455 -41 461 -36
rect 466 -39 478 -35
rect 482 -39 483 -35
rect 487 -39 488 -35
rect 455 -43 457 -41
rect 448 -45 457 -43
rect 487 -40 492 -39
rect 496 -39 500 -23
rect 524 -20 529 -17
rect 524 -24 525 -20
rect 550 -20 561 -16
rect 550 -24 554 -20
rect 568 -23 569 -19
rect 573 -23 584 -19
rect 524 -25 529 -24
rect 533 -26 554 -24
rect 525 -30 533 -29
rect 537 -28 554 -26
rect 525 -33 537 -30
rect 487 -44 491 -40
rect 448 -49 461 -45
rect 467 -48 491 -44
rect 496 -43 498 -39
rect 441 -50 445 -49
rect 467 -50 471 -48
rect 454 -57 455 -53
rect 459 -57 460 -53
rect 496 -52 500 -43
rect 525 -45 529 -33
rect 550 -35 554 -28
rect 558 -30 559 -26
rect 563 -27 564 -26
rect 563 -30 575 -27
rect 558 -31 575 -30
rect 571 -34 575 -31
rect 571 -35 576 -34
rect 539 -41 545 -36
rect 550 -39 562 -35
rect 566 -39 567 -35
rect 571 -39 572 -35
rect 539 -43 541 -41
rect 532 -45 541 -43
rect 571 -40 576 -39
rect 571 -44 575 -40
rect 532 -49 545 -45
rect 551 -48 575 -44
rect 525 -50 529 -49
rect 551 -50 555 -48
rect 467 -55 471 -54
rect 476 -56 477 -52
rect 481 -56 500 -52
rect 454 -62 460 -57
rect 538 -57 539 -53
rect 543 -57 544 -53
rect 580 -52 584 -23
rect 594 -26 598 -19
rect 594 -27 599 -26
rect 594 -31 595 -27
rect 602 -27 606 -6
rect 609 -12 622 -11
rect 609 -16 612 -12
rect 616 -16 618 -12
rect 609 -17 622 -16
rect 609 -24 615 -17
rect 625 -23 629 -6
rect 602 -31 605 -27
rect 609 -31 610 -27
rect 614 -31 615 -27
rect 619 -31 620 -27
rect 625 -28 629 -27
rect 594 -32 599 -31
rect 594 -40 598 -32
rect 614 -36 620 -31
rect 601 -40 602 -36
rect 606 -40 620 -36
rect 626 -37 630 -35
rect 551 -55 555 -54
rect 560 -56 561 -52
rect 565 -56 584 -52
rect 588 -43 598 -40
rect 588 -55 591 -43
rect 538 -62 544 -57
rect 594 -49 598 -43
rect 594 -50 599 -49
rect 594 -54 595 -50
rect 599 -54 606 -51
rect 594 -57 606 -54
rect 610 -53 614 -40
rect 626 -44 630 -41
rect 617 -48 621 -44
rect 625 -48 630 -44
rect 617 -49 630 -48
rect 610 -57 624 -53
rect 628 -57 629 -53
rect 361 -66 364 -62
rect 368 -66 374 -62
rect 378 -66 442 -62
rect 446 -66 495 -62
rect 499 -66 526 -62
rect 530 -66 579 -62
rect 583 -66 596 -62
rect 600 -66 606 -62
rect 610 -66 634 -62
rect 342 -69 627 -66
rect 361 -70 627 -69
rect 631 -70 634 -66
rect 451 -72 495 -70
rect 451 -76 457 -72
rect 461 -76 485 -72
rect 489 -76 495 -72
rect 422 -81 425 -79
rect 455 -84 461 -76
rect 422 -99 425 -85
rect 455 -88 456 -84
rect 460 -88 461 -84
rect 466 -84 470 -83
rect 475 -84 481 -76
rect 475 -88 476 -84
rect 480 -88 481 -84
rect 486 -84 491 -81
rect 490 -88 491 -84
rect 466 -91 470 -88
rect 486 -89 491 -88
rect 466 -95 483 -91
rect 327 -137 332 -117
rect 394 -103 422 -100
rect 394 -129 398 -103
rect 455 -107 459 -97
rect 463 -102 468 -98
rect 479 -99 483 -95
rect 463 -110 469 -106
rect 473 -110 476 -106
rect 463 -116 467 -110
rect 479 -114 483 -103
rect 450 -119 467 -116
rect 471 -118 483 -114
rect 471 -122 475 -118
rect 487 -119 491 -89
rect 518 -93 600 -88
rect 655 -114 659 -3
rect 689 -23 693 -16
rect 689 -24 694 -23
rect 689 -28 690 -24
rect 697 -24 701 -3
rect 704 -9 717 -8
rect 704 -13 707 -9
rect 711 -13 713 -9
rect 704 -14 717 -13
rect 704 -21 710 -14
rect 720 -20 724 -3
rect 790 -3 802 -2
rect 806 -2 886 1
rect 806 -3 870 -2
rect 767 -14 779 -8
rect 786 -9 790 -6
rect 874 -3 886 -2
rect 890 -3 923 1
rect 927 -3 937 1
rect 941 -3 951 1
rect 955 -3 961 1
rect 800 -12 822 -8
rect 826 -12 827 -8
rect 851 -9 863 -8
rect 800 -13 804 -12
rect 786 -14 790 -13
rect 767 -17 772 -14
rect 767 -18 768 -17
rect 697 -28 700 -24
rect 704 -28 705 -24
rect 709 -28 710 -24
rect 714 -28 715 -24
rect 720 -25 724 -24
rect 759 -21 768 -18
rect 793 -17 804 -13
rect 851 -13 856 -9
rect 860 -13 863 -9
rect 851 -14 863 -13
rect 870 -9 874 -6
rect 884 -12 906 -8
rect 910 -12 911 -8
rect 884 -13 888 -12
rect 870 -14 874 -13
rect 793 -21 797 -17
rect 811 -20 812 -16
rect 816 -20 827 -16
rect 689 -29 694 -28
rect 689 -37 693 -29
rect 709 -33 715 -28
rect 696 -37 697 -33
rect 701 -37 715 -33
rect 721 -35 725 -32
rect 759 -35 762 -21
rect 767 -22 772 -21
rect 776 -23 797 -21
rect 689 -46 693 -41
rect 689 -47 694 -46
rect 689 -51 690 -47
rect 694 -51 701 -48
rect 689 -54 701 -51
rect 705 -50 709 -37
rect 768 -27 776 -26
rect 780 -25 797 -23
rect 768 -30 780 -27
rect 721 -41 725 -39
rect 712 -45 716 -41
rect 720 -45 725 -41
rect 712 -46 725 -45
rect 768 -42 772 -30
rect 793 -32 797 -25
rect 801 -27 802 -23
rect 806 -24 807 -23
rect 806 -27 818 -24
rect 801 -28 818 -27
rect 814 -31 818 -28
rect 814 -32 819 -31
rect 782 -38 788 -33
rect 793 -36 805 -32
rect 809 -36 810 -32
rect 814 -36 815 -32
rect 782 -40 784 -38
rect 768 -47 772 -46
rect 775 -42 784 -40
rect 814 -37 819 -36
rect 823 -36 827 -20
rect 851 -17 856 -14
rect 851 -21 852 -17
rect 877 -17 888 -13
rect 877 -21 881 -17
rect 895 -20 896 -16
rect 900 -20 911 -16
rect 851 -22 856 -21
rect 860 -23 881 -21
rect 852 -27 860 -26
rect 864 -25 881 -23
rect 852 -30 864 -27
rect 814 -41 818 -37
rect 775 -46 788 -42
rect 794 -45 818 -41
rect 823 -40 825 -36
rect 705 -54 719 -50
rect 723 -54 724 -50
rect 775 -51 778 -46
rect 794 -47 798 -45
rect 764 -55 778 -51
rect 781 -54 782 -50
rect 786 -54 787 -50
rect 823 -49 827 -40
rect 852 -42 856 -30
rect 877 -32 881 -25
rect 885 -27 886 -23
rect 890 -24 891 -23
rect 890 -27 902 -24
rect 885 -28 902 -27
rect 898 -31 902 -28
rect 898 -32 903 -31
rect 866 -38 872 -33
rect 877 -36 889 -32
rect 893 -36 894 -32
rect 898 -36 899 -32
rect 866 -40 868 -38
rect 859 -42 868 -40
rect 898 -37 903 -36
rect 898 -41 902 -37
rect 859 -46 872 -42
rect 878 -45 902 -41
rect 852 -47 856 -46
rect 878 -47 882 -45
rect 794 -52 798 -51
rect 803 -53 804 -49
rect 808 -53 827 -49
rect 764 -59 768 -55
rect 781 -59 787 -54
rect 865 -54 866 -50
rect 870 -54 871 -50
rect 907 -49 911 -20
rect 921 -23 925 -16
rect 921 -24 926 -23
rect 921 -28 922 -24
rect 929 -24 933 -3
rect 936 -9 949 -8
rect 936 -13 939 -9
rect 943 -13 945 -9
rect 936 -14 949 -13
rect 936 -21 942 -14
rect 952 -20 956 -3
rect 929 -28 932 -24
rect 936 -28 937 -24
rect 941 -28 942 -24
rect 946 -28 947 -24
rect 952 -25 956 -24
rect 921 -29 926 -28
rect 921 -37 925 -29
rect 941 -33 947 -28
rect 928 -37 929 -33
rect 933 -37 947 -33
rect 953 -34 957 -32
rect 878 -52 882 -51
rect 887 -53 888 -49
rect 892 -53 911 -49
rect 915 -40 925 -37
rect 915 -52 918 -40
rect 865 -59 871 -54
rect 921 -46 925 -40
rect 921 -47 926 -46
rect 921 -51 922 -47
rect 926 -51 933 -48
rect 921 -54 933 -51
rect 937 -50 941 -37
rect 953 -41 957 -38
rect 944 -45 948 -41
rect 952 -45 957 -41
rect 944 -46 957 -45
rect 937 -54 951 -50
rect 955 -54 956 -50
rect 688 -62 691 -59
rect 687 -63 691 -62
rect 695 -63 701 -59
rect 705 -63 769 -59
rect 773 -63 822 -59
rect 826 -63 853 -59
rect 857 -63 906 -59
rect 910 -63 923 -59
rect 927 -63 933 -59
rect 937 -63 961 -59
rect 687 -65 961 -63
rect 668 -66 961 -65
rect 671 -67 961 -66
rect 671 -68 690 -67
rect 778 -69 822 -67
rect 778 -73 784 -69
rect 788 -73 812 -69
rect 816 -73 822 -69
rect 725 -75 729 -74
rect 669 -93 698 -88
rect 486 -120 491 -119
rect 455 -126 456 -122
rect 460 -126 475 -122
rect 478 -124 486 -122
rect 490 -122 491 -120
rect 490 -124 495 -122
rect 478 -126 495 -124
rect 473 -132 474 -129
rect 451 -133 474 -132
rect 478 -132 479 -129
rect 478 -133 485 -132
rect 451 -136 485 -133
rect 489 -136 495 -132
rect 451 -137 495 -136
rect 327 -140 495 -137
rect 654 -134 659 -114
rect 725 -116 729 -79
rect 782 -81 788 -73
rect 782 -85 783 -81
rect 787 -85 788 -81
rect 793 -81 797 -80
rect 802 -81 808 -73
rect 802 -85 803 -81
rect 807 -85 808 -81
rect 813 -81 818 -78
rect 817 -85 818 -81
rect 793 -88 797 -85
rect 813 -86 818 -85
rect 793 -92 810 -88
rect 782 -104 786 -94
rect 790 -99 795 -95
rect 806 -96 810 -92
rect 790 -107 796 -103
rect 800 -107 803 -103
rect 790 -113 794 -107
rect 806 -111 810 -100
rect 777 -116 794 -113
rect 798 -115 810 -111
rect 814 -91 830 -86
rect 798 -119 802 -115
rect 814 -116 818 -91
rect 813 -117 818 -116
rect 782 -123 783 -119
rect 787 -123 802 -119
rect 805 -121 813 -119
rect 817 -121 818 -117
rect 805 -123 818 -121
rect 800 -129 801 -126
rect 778 -130 801 -129
rect 805 -129 806 -126
rect 805 -130 812 -129
rect 778 -133 812 -130
rect 816 -133 822 -129
rect 778 -134 822 -133
rect 654 -137 822 -134
rect 654 -138 778 -137
rect 327 -141 451 -140
rect 440 -148 444 -141
rect 323 -150 367 -148
rect 416 -150 460 -148
rect 503 -150 547 -148
rect 323 -152 547 -150
rect 323 -156 329 -152
rect 333 -153 422 -152
rect 333 -156 367 -153
rect 416 -156 422 -153
rect 426 -153 509 -152
rect 426 -156 460 -153
rect 503 -156 509 -153
rect 513 -156 547 -152
rect 337 -164 343 -156
rect 337 -168 338 -164
rect 342 -168 343 -164
rect 348 -162 352 -161
rect 357 -162 363 -156
rect 398 -162 409 -159
rect 357 -166 358 -162
rect 362 -166 363 -162
rect 327 -169 332 -168
rect 327 -173 328 -169
rect 348 -169 352 -166
rect 327 -176 332 -173
rect 327 -180 328 -176
rect 327 -181 332 -180
rect 335 -173 348 -171
rect 335 -175 352 -173
rect 359 -173 390 -169
rect 327 -182 331 -181
rect 291 -186 331 -182
rect 327 -199 331 -186
rect 335 -186 339 -175
rect 350 -182 355 -178
rect 359 -182 363 -173
rect 342 -190 345 -186
rect 349 -190 356 -186
rect 335 -194 339 -190
rect 335 -198 347 -194
rect 351 -195 356 -190
rect 327 -200 332 -199
rect 327 -204 328 -200
rect 332 -204 339 -201
rect 327 -207 339 -204
rect 343 -202 347 -198
rect 350 -199 366 -195
rect 343 -206 358 -202
rect 362 -206 363 -202
rect 386 -206 390 -173
rect 406 -172 409 -162
rect 430 -164 436 -156
rect 430 -168 431 -164
rect 435 -168 436 -164
rect 441 -162 445 -161
rect 450 -162 456 -156
rect 450 -166 451 -162
rect 455 -166 456 -162
rect 517 -164 523 -156
rect 496 -165 512 -164
rect 420 -169 425 -168
rect 420 -172 421 -169
rect 406 -173 421 -172
rect 441 -169 445 -166
rect 406 -175 425 -173
rect 420 -176 425 -175
rect 420 -180 421 -176
rect 420 -181 425 -180
rect 428 -173 441 -171
rect 428 -175 445 -173
rect 420 -199 424 -181
rect 428 -186 432 -175
rect 452 -178 456 -169
rect 500 -169 512 -165
rect 517 -168 518 -164
rect 522 -168 523 -164
rect 528 -162 532 -161
rect 537 -162 543 -156
rect 537 -166 538 -162
rect 542 -166 543 -162
rect 500 -170 508 -169
rect 507 -173 508 -170
rect 528 -169 532 -166
rect 507 -176 512 -173
rect 443 -182 448 -178
rect 452 -182 463 -178
rect 507 -180 508 -176
rect 507 -181 512 -180
rect 515 -173 528 -171
rect 515 -175 532 -173
rect 435 -190 438 -186
rect 442 -190 449 -186
rect 428 -194 432 -190
rect 428 -198 440 -194
rect 420 -200 425 -199
rect 420 -204 421 -200
rect 425 -204 432 -201
rect 420 -207 432 -204
rect 436 -202 440 -198
rect 444 -195 449 -190
rect 444 -199 459 -195
rect 507 -199 511 -181
rect 515 -186 519 -175
rect 539 -178 543 -169
rect 530 -182 535 -178
rect 539 -182 552 -178
rect 522 -190 525 -186
rect 529 -190 536 -186
rect 515 -194 519 -190
rect 515 -198 527 -194
rect 507 -200 512 -199
rect 436 -206 451 -202
rect 455 -206 456 -202
rect 507 -204 508 -200
rect 512 -204 519 -201
rect 507 -207 519 -204
rect 523 -202 527 -198
rect 531 -196 536 -190
rect 531 -199 544 -196
rect 523 -206 538 -202
rect 542 -206 543 -202
rect 323 -216 329 -212
rect 333 -216 339 -212
rect 343 -216 367 -212
rect 416 -216 422 -212
rect 426 -216 432 -212
rect 436 -216 460 -212
rect 317 -217 460 -216
rect 503 -216 509 -212
rect 513 -216 519 -212
rect 523 -216 547 -212
rect 503 -217 547 -216
rect 317 -219 547 -217
rect 323 -220 367 -219
rect 416 -220 547 -219
<< metal2 >>
rect 79 224 108 228
rect 15 220 82 224
rect 15 78 20 220
rect 89 213 342 217
rect 30 155 34 206
rect 89 178 94 213
rect 337 209 341 213
rect 107 200 108 203
rect 112 200 196 203
rect 200 200 289 203
rect 472 199 476 233
rect 514 214 762 218
rect 514 210 518 214
rect 571 202 660 205
rect 569 201 660 202
rect 664 201 747 205
rect 193 182 337 185
rect 519 184 666 187
rect 88 174 100 178
rect 193 178 196 182
rect 663 180 666 184
rect 105 174 116 178
rect 245 173 246 176
rect 29 153 34 155
rect 29 117 33 153
rect 173 152 221 155
rect 173 151 230 152
rect 218 148 230 151
rect 243 142 246 173
rect 286 168 289 174
rect 567 176 571 179
rect 286 165 337 168
rect 567 168 570 176
rect 519 165 570 168
rect 663 176 664 180
rect 681 178 700 182
rect 758 180 762 214
rect 744 176 752 180
rect 757 178 762 180
rect 757 176 984 178
rect 564 157 567 165
rect 491 154 502 156
rect 564 154 578 157
rect 491 153 496 154
rect 272 150 496 153
rect 500 150 502 154
rect 272 149 502 150
rect 602 148 605 175
rect 664 166 667 176
rect 758 175 984 176
rect 771 174 984 175
rect 970 166 974 167
rect 664 162 974 166
rect 617 154 676 157
rect 507 145 605 148
rect 704 154 966 157
rect 690 150 694 153
rect 690 147 757 150
rect 195 141 248 142
rect 113 138 248 141
rect 507 140 511 145
rect 113 132 116 138
rect 62 129 127 132
rect 29 113 70 117
rect 66 106 70 113
rect 19 74 20 78
rect 27 104 30 105
rect 27 101 34 104
rect 27 36 30 101
rect 70 102 103 105
rect 123 105 126 129
rect 205 129 290 132
rect 294 129 315 132
rect 391 131 456 134
rect 174 101 207 104
rect 187 97 190 101
rect 299 97 302 103
rect 187 94 302 97
rect 263 85 264 88
rect 261 37 264 85
rect 312 79 315 129
rect 452 128 456 131
rect 507 128 510 140
rect 753 137 757 147
rect 514 134 534 136
rect 514 133 530 134
rect 514 129 515 133
rect 519 130 530 133
rect 534 131 619 134
rect 718 134 783 137
rect 519 129 534 130
rect 514 128 522 129
rect 452 125 510 128
rect 356 103 363 106
rect 306 75 340 79
rect 300 74 340 75
rect 27 33 121 36
rect 131 34 274 37
rect 118 29 121 33
rect 269 3 300 7
rect 250 2 274 3
rect 207 -1 274 2
rect 207 -2 210 -1
rect 151 -5 210 -2
rect 151 -14 155 -5
rect 61 -17 155 -14
rect 26 -45 33 -42
rect 26 -110 29 -45
rect 69 -44 102 -41
rect 122 -41 125 -17
rect 204 -17 289 -14
rect 83 -79 86 -44
rect 173 -45 206 -42
rect 186 -49 189 -45
rect 298 -49 301 -43
rect 186 -52 301 -49
rect 262 -61 263 -58
rect 183 -77 186 -61
rect 83 -83 176 -79
rect 182 -80 249 -77
rect 171 -96 176 -83
rect 171 -100 244 -96
rect 260 -109 263 -61
rect 313 -65 316 74
rect 324 51 345 55
rect 356 38 359 103
rect 399 104 432 107
rect 452 107 455 125
rect 591 123 749 126
rect 417 55 421 104
rect 503 103 536 106
rect 516 99 519 103
rect 628 99 631 105
rect 516 96 631 99
rect 683 106 690 109
rect 592 87 593 90
rect 590 39 593 87
rect 633 77 667 81
rect 627 76 667 77
rect 643 48 671 51
rect 683 41 686 106
rect 726 107 759 110
rect 779 110 782 134
rect 861 134 946 137
rect 838 126 912 128
rect 838 125 916 126
rect 742 52 746 107
rect 830 106 863 109
rect 843 102 846 106
rect 955 102 958 108
rect 843 99 958 102
rect 751 65 754 90
rect 919 90 920 93
rect 768 53 827 56
rect 835 52 839 90
rect 917 42 920 90
rect 356 35 450 38
rect 460 36 603 39
rect 683 38 777 41
rect 787 39 930 42
rect 447 31 450 35
rect 774 34 777 38
rect 745 27 765 30
rect 745 25 748 27
rect 505 22 748 25
rect 762 26 765 27
rect 825 27 873 30
rect 762 22 764 26
rect 768 22 769 25
rect 505 6 508 22
rect 825 18 828 27
rect 756 16 828 18
rect 752 15 828 16
rect 834 9 839 12
rect 325 3 508 6
rect 534 5 839 9
rect 534 4 657 5
rect 535 -12 540 4
rect 867 -9 870 27
rect 390 -15 455 -12
rect 422 -31 425 -15
rect 355 -43 362 -40
rect 308 -66 338 -65
rect 308 -71 337 -66
rect 278 -100 298 -96
rect 26 -113 120 -110
rect 130 -112 273 -109
rect 117 -117 120 -113
rect 309 -214 315 -71
rect 336 -96 340 -95
rect 324 -100 340 -96
rect 336 -121 340 -100
rect 355 -108 358 -43
rect 398 -42 431 -39
rect 451 -39 454 -15
rect 533 -15 618 -12
rect 717 -12 782 -9
rect 413 -89 416 -42
rect 502 -43 535 -40
rect 515 -47 518 -43
rect 627 -47 630 -41
rect 515 -50 630 -47
rect 682 -40 689 -37
rect 422 -55 425 -54
rect 591 -59 592 -56
rect 422 -81 425 -59
rect 413 -93 512 -89
rect 589 -107 592 -59
rect 631 -69 667 -66
rect 605 -93 664 -88
rect 682 -105 685 -40
rect 725 -39 758 -36
rect 778 -36 781 -12
rect 860 -12 945 -9
rect 745 -75 749 -39
rect 829 -40 862 -37
rect 842 -44 845 -40
rect 954 -44 957 -38
rect 842 -47 957 -44
rect 918 -56 919 -53
rect 729 -79 749 -75
rect 745 -80 749 -79
rect 703 -91 830 -88
rect 836 -91 837 -88
rect 703 -92 837 -91
rect 916 -104 919 -56
rect 355 -111 449 -108
rect 459 -110 602 -107
rect 682 -108 776 -105
rect 786 -107 929 -104
rect 446 -115 449 -111
rect 773 -112 776 -108
rect 725 -116 729 -115
rect 336 -125 413 -121
rect 410 -129 413 -125
rect 493 -126 495 -121
rect 493 -129 498 -126
rect 394 -158 398 -133
rect 410 -133 498 -129
rect 410 -134 413 -133
rect 725 -165 729 -120
rect 963 -126 966 154
rect 500 -168 729 -165
rect 500 -169 725 -168
rect 962 -178 966 -126
rect 467 -182 501 -178
rect 556 -181 966 -178
rect 962 -182 966 -181
rect 497 -186 501 -182
rect 497 -189 566 -186
rect 563 -193 566 -189
rect 970 -193 974 162
rect 371 -199 459 -195
rect 464 -199 544 -196
rect 563 -197 974 -193
rect 981 -207 984 174
rect 390 -210 984 -207
rect 309 -221 310 -214
<< metal3 >>
rect 495 154 520 156
rect 495 150 496 154
rect 500 150 520 154
rect 495 149 501 150
rect 514 135 520 150
rect 514 133 521 135
rect 514 129 515 133
rect 519 129 521 133
rect 514 128 521 129
<< ntransistor >>
rect 119 201 121 212
rect 126 201 128 212
rect 139 201 141 210
rect 206 201 208 212
rect 213 201 215 212
rect 226 201 228 210
rect 299 201 301 212
rect 306 201 308 212
rect 319 201 321 210
rect 539 203 541 212
rect 552 203 554 214
rect 559 203 561 214
rect 632 203 634 212
rect 645 203 647 214
rect 652 203 654 214
rect 719 203 721 212
rect 732 203 734 214
rect 739 203 741 214
rect 41 89 43 95
rect 53 83 55 92
rect 60 83 62 92
rect 119 91 121 100
rect 135 86 137 95
rect 145 86 147 95
rect 155 83 157 95
rect 162 83 164 95
rect 203 91 205 100
rect 219 86 221 95
rect 229 86 231 95
rect 239 83 241 95
rect 246 83 248 95
rect 273 89 275 95
rect 285 83 287 92
rect 292 83 294 92
rect 370 91 372 97
rect 382 85 384 94
rect 389 85 391 94
rect 448 93 450 102
rect 464 88 466 97
rect 474 88 476 97
rect 484 85 486 97
rect 491 85 493 97
rect 532 93 534 102
rect 548 88 550 97
rect 558 88 560 97
rect 568 85 570 97
rect 575 85 577 97
rect 602 91 604 97
rect 697 94 699 100
rect 614 85 616 94
rect 621 85 623 94
rect 709 88 711 97
rect 716 88 718 97
rect 775 96 777 105
rect 791 91 793 100
rect 801 91 803 100
rect 811 88 813 100
rect 818 88 820 100
rect 859 96 861 105
rect 875 91 877 100
rect 885 91 887 100
rect 895 88 897 100
rect 902 88 904 100
rect 929 94 931 100
rect 941 88 943 97
rect 948 88 950 97
rect 134 55 136 61
rect 144 55 146 61
rect 154 55 156 61
rect 463 57 465 63
rect 473 57 475 63
rect 483 57 485 63
rect 790 60 792 66
rect 800 60 802 66
rect 810 60 812 66
rect 40 -57 42 -51
rect 52 -63 54 -54
rect 59 -63 61 -54
rect 118 -55 120 -46
rect 134 -60 136 -51
rect 144 -60 146 -51
rect 154 -63 156 -51
rect 161 -63 163 -51
rect 202 -55 204 -46
rect 218 -60 220 -51
rect 228 -60 230 -51
rect 238 -63 240 -51
rect 245 -63 247 -51
rect 272 -57 274 -51
rect 284 -63 286 -54
rect 291 -63 293 -54
rect 369 -55 371 -49
rect 381 -61 383 -52
rect 388 -61 390 -52
rect 447 -53 449 -44
rect 463 -58 465 -49
rect 473 -58 475 -49
rect 483 -61 485 -49
rect 490 -61 492 -49
rect 531 -53 533 -44
rect 547 -58 549 -49
rect 557 -58 559 -49
rect 567 -61 569 -49
rect 574 -61 576 -49
rect 601 -55 603 -49
rect 696 -52 698 -46
rect 613 -61 615 -52
rect 620 -61 622 -52
rect 708 -58 710 -49
rect 715 -58 717 -49
rect 774 -50 776 -41
rect 790 -55 792 -46
rect 800 -55 802 -46
rect 810 -58 812 -46
rect 817 -58 819 -46
rect 858 -50 860 -41
rect 874 -55 876 -46
rect 884 -55 886 -46
rect 894 -58 896 -46
rect 901 -58 903 -46
rect 928 -52 930 -46
rect 940 -58 942 -49
rect 947 -58 949 -49
rect 133 -91 135 -85
rect 143 -91 145 -85
rect 153 -91 155 -85
rect 462 -89 464 -83
rect 472 -89 474 -83
rect 482 -89 484 -83
rect 789 -86 791 -80
rect 799 -86 801 -80
rect 809 -86 811 -80
rect 334 -205 336 -196
rect 347 -207 349 -196
rect 354 -207 356 -196
rect 427 -205 429 -196
rect 440 -207 442 -196
rect 447 -207 449 -196
rect 514 -205 516 -196
rect 527 -207 529 -196
rect 534 -207 536 -196
<< ptransistor >>
rect 119 166 121 179
rect 129 166 131 179
rect 139 168 141 186
rect 206 166 208 179
rect 216 166 218 179
rect 226 168 228 186
rect 299 166 301 179
rect 309 166 311 179
rect 319 168 321 186
rect 539 170 541 188
rect 549 168 551 181
rect 559 168 561 181
rect 632 170 634 188
rect 642 168 644 181
rect 652 168 654 181
rect 719 170 721 188
rect 729 168 731 181
rect 739 168 741 181
rect 41 112 43 124
rect 51 112 53 122
rect 61 112 63 122
rect 127 113 129 140
rect 143 113 145 131
rect 153 113 155 131
rect 163 113 165 140
rect 211 113 213 140
rect 227 113 229 131
rect 237 113 239 131
rect 247 113 249 140
rect 273 112 275 124
rect 283 112 285 122
rect 293 112 295 122
rect 370 114 372 126
rect 380 114 382 124
rect 390 114 392 124
rect 456 115 458 142
rect 472 115 474 133
rect 482 115 484 133
rect 492 115 494 142
rect 540 115 542 142
rect 556 115 558 133
rect 566 115 568 133
rect 576 115 578 142
rect 602 114 604 126
rect 612 114 614 124
rect 622 114 624 124
rect 697 117 699 129
rect 707 117 709 127
rect 717 117 719 127
rect 783 118 785 145
rect 799 118 801 136
rect 809 118 811 136
rect 819 118 821 145
rect 867 118 869 145
rect 883 118 885 136
rect 893 118 895 136
rect 903 118 905 145
rect 929 117 931 129
rect 939 117 941 127
rect 949 117 951 127
rect 134 10 136 28
rect 141 10 143 28
rect 154 19 156 31
rect 463 12 465 30
rect 470 12 472 30
rect 483 21 485 33
rect 790 15 792 33
rect 797 15 799 33
rect 810 24 812 36
rect 40 -34 42 -22
rect 50 -34 52 -24
rect 60 -34 62 -24
rect 126 -33 128 -6
rect 142 -33 144 -15
rect 152 -33 154 -15
rect 162 -33 164 -6
rect 210 -33 212 -6
rect 226 -33 228 -15
rect 236 -33 238 -15
rect 246 -33 248 -6
rect 272 -34 274 -22
rect 282 -34 284 -24
rect 292 -34 294 -24
rect 369 -32 371 -20
rect 379 -32 381 -22
rect 389 -32 391 -22
rect 455 -31 457 -4
rect 471 -31 473 -13
rect 481 -31 483 -13
rect 491 -31 493 -4
rect 539 -31 541 -4
rect 555 -31 557 -13
rect 565 -31 567 -13
rect 575 -31 577 -4
rect 601 -32 603 -20
rect 611 -32 613 -22
rect 621 -32 623 -22
rect 696 -29 698 -17
rect 706 -29 708 -19
rect 716 -29 718 -19
rect 782 -28 784 -1
rect 798 -28 800 -10
rect 808 -28 810 -10
rect 818 -28 820 -1
rect 866 -28 868 -1
rect 882 -28 884 -10
rect 892 -28 894 -10
rect 902 -28 904 -1
rect 928 -29 930 -17
rect 938 -29 940 -19
rect 948 -29 950 -19
rect 133 -136 135 -118
rect 140 -136 142 -118
rect 153 -127 155 -115
rect 462 -134 464 -116
rect 469 -134 471 -116
rect 482 -125 484 -113
rect 789 -131 791 -113
rect 796 -131 798 -113
rect 809 -122 811 -110
rect 334 -181 336 -163
rect 344 -174 346 -161
rect 354 -174 356 -161
rect 427 -181 429 -163
rect 437 -174 439 -161
rect 447 -174 449 -161
rect 514 -181 516 -163
rect 524 -174 526 -161
rect 534 -174 536 -161
<< polycontact >>
rect 126 191 130 195
rect 136 191 140 195
rect 116 183 120 187
rect 213 191 217 195
rect 223 191 227 195
rect 203 183 207 187
rect 306 191 310 195
rect 316 191 320 195
rect 296 183 300 187
rect 540 193 544 197
rect 550 193 554 197
rect 633 193 637 197
rect 643 193 647 197
rect 560 185 564 189
rect 720 193 724 197
rect 730 193 734 197
rect 653 185 657 189
rect 740 185 744 189
rect 52 128 56 132
rect 113 120 117 124
rect 42 104 46 108
rect 197 120 201 124
rect 150 105 154 109
rect 160 105 164 109
rect 284 128 288 132
rect 381 130 385 134
rect 442 122 446 126
rect 61 96 65 100
rect 129 99 133 103
rect 234 105 238 109
rect 244 105 248 109
rect 274 104 278 108
rect 213 99 217 103
rect 371 106 375 110
rect 293 96 297 100
rect 526 122 530 126
rect 479 107 483 111
rect 489 107 493 111
rect 613 130 617 134
rect 708 133 712 137
rect 769 125 773 129
rect 390 98 394 102
rect 458 101 462 105
rect 563 107 567 111
rect 573 107 577 111
rect 603 106 607 110
rect 542 101 546 105
rect 698 109 702 113
rect 622 98 626 102
rect 853 125 857 129
rect 806 110 810 114
rect 816 110 820 114
rect 940 133 944 137
rect 717 101 721 105
rect 785 104 789 108
rect 890 110 894 114
rect 900 110 904 114
rect 930 109 934 113
rect 869 104 873 108
rect 949 101 953 105
rect 131 42 135 46
rect 143 42 147 46
rect 151 41 155 45
rect 460 44 464 48
rect 472 44 476 48
rect 141 34 145 38
rect 480 43 484 47
rect 787 47 791 51
rect 799 47 803 51
rect 470 36 474 40
rect 807 46 811 50
rect 797 39 801 43
rect 51 -18 55 -14
rect 112 -26 116 -22
rect 41 -42 45 -38
rect 196 -26 200 -22
rect 149 -41 153 -37
rect 159 -41 163 -37
rect 283 -18 287 -14
rect 380 -16 384 -12
rect 441 -24 445 -20
rect 60 -50 64 -46
rect 128 -47 132 -43
rect 233 -41 237 -37
rect 243 -41 247 -37
rect 273 -42 277 -38
rect 212 -47 216 -43
rect 370 -40 374 -36
rect 292 -50 296 -46
rect 525 -24 529 -20
rect 478 -39 482 -35
rect 488 -39 492 -35
rect 612 -16 616 -12
rect 707 -13 711 -9
rect 768 -21 772 -17
rect 389 -48 393 -44
rect 457 -45 461 -41
rect 562 -39 566 -35
rect 572 -39 576 -35
rect 602 -40 606 -36
rect 541 -45 545 -41
rect 697 -37 701 -33
rect 621 -48 625 -44
rect 852 -21 856 -17
rect 805 -36 809 -32
rect 815 -36 819 -32
rect 939 -13 943 -9
rect 716 -45 720 -41
rect 784 -42 788 -38
rect 889 -36 893 -32
rect 899 -36 903 -32
rect 929 -37 933 -33
rect 868 -42 872 -38
rect 948 -45 952 -41
rect 130 -104 134 -100
rect 142 -104 146 -100
rect 150 -105 154 -101
rect 459 -102 463 -98
rect 471 -102 475 -98
rect 140 -112 144 -108
rect 479 -103 483 -99
rect 786 -99 790 -95
rect 798 -99 802 -95
rect 469 -110 473 -106
rect 806 -100 810 -96
rect 796 -107 800 -103
rect 355 -182 359 -178
rect 335 -190 339 -186
rect 345 -190 349 -186
rect 448 -182 452 -178
rect 428 -190 432 -186
rect 438 -190 442 -186
rect 535 -182 539 -178
rect 515 -190 519 -186
rect 525 -190 529 -186
<< ndcontact >>
rect 132 217 136 221
rect 219 217 223 221
rect 113 207 117 211
rect 312 217 316 221
rect 143 205 147 209
rect 200 207 204 211
rect 544 219 548 223
rect 230 205 234 209
rect 293 207 297 211
rect 637 219 641 223
rect 323 205 327 209
rect 533 207 537 211
rect 563 209 567 213
rect 724 219 728 223
rect 626 207 630 211
rect 656 209 660 213
rect 713 207 717 211
rect 743 209 747 213
rect 35 90 39 94
rect 113 95 117 99
rect 197 95 201 99
rect 64 87 68 91
rect 127 87 131 91
rect 139 90 143 94
rect 149 88 153 92
rect 46 78 50 82
rect 211 87 215 91
rect 223 90 227 94
rect 233 88 237 92
rect 167 78 171 82
rect 267 90 271 94
rect 364 92 368 96
rect 442 97 446 101
rect 296 87 300 91
rect 526 97 530 101
rect 393 89 397 93
rect 456 89 460 93
rect 468 92 472 96
rect 478 90 482 94
rect 251 78 255 82
rect 278 78 282 82
rect 375 80 379 84
rect 540 89 544 93
rect 552 92 556 96
rect 562 90 566 94
rect 496 80 500 84
rect 596 92 600 96
rect 691 95 695 99
rect 769 100 773 104
rect 625 89 629 93
rect 853 100 857 104
rect 720 92 724 96
rect 783 92 787 96
rect 795 95 799 99
rect 805 93 809 97
rect 580 80 584 84
rect 607 80 611 84
rect 702 83 706 87
rect 867 92 871 96
rect 879 95 883 99
rect 889 93 893 97
rect 823 83 827 87
rect 923 95 927 99
rect 952 92 956 96
rect 907 83 911 87
rect 934 83 938 87
rect 128 56 132 60
rect 138 56 142 60
rect 148 56 152 60
rect 158 56 162 60
rect 457 58 461 62
rect 467 58 471 62
rect 477 58 481 62
rect 487 58 491 62
rect 784 61 788 65
rect 794 61 798 65
rect 804 61 808 65
rect 814 61 818 65
rect 34 -56 38 -52
rect 112 -51 116 -47
rect 196 -51 200 -47
rect 63 -59 67 -55
rect 126 -59 130 -55
rect 138 -56 142 -52
rect 148 -58 152 -54
rect 45 -68 49 -64
rect 210 -59 214 -55
rect 222 -56 226 -52
rect 232 -58 236 -54
rect 166 -68 170 -64
rect 266 -56 270 -52
rect 363 -54 367 -50
rect 441 -49 445 -45
rect 295 -59 299 -55
rect 525 -49 529 -45
rect 392 -57 396 -53
rect 455 -57 459 -53
rect 467 -54 471 -50
rect 477 -56 481 -52
rect 250 -68 254 -64
rect 277 -68 281 -64
rect 374 -66 378 -62
rect 539 -57 543 -53
rect 551 -54 555 -50
rect 561 -56 565 -52
rect 495 -66 499 -62
rect 595 -54 599 -50
rect 690 -51 694 -47
rect 768 -46 772 -42
rect 624 -57 628 -53
rect 852 -46 856 -42
rect 719 -54 723 -50
rect 782 -54 786 -50
rect 794 -51 798 -47
rect 804 -53 808 -49
rect 579 -66 583 -62
rect 606 -66 610 -62
rect 701 -63 705 -59
rect 866 -54 870 -50
rect 878 -51 882 -47
rect 888 -53 892 -49
rect 822 -63 826 -59
rect 922 -51 926 -47
rect 951 -54 955 -50
rect 906 -63 910 -59
rect 933 -63 937 -59
rect 127 -90 131 -86
rect 137 -90 141 -86
rect 147 -90 151 -86
rect 157 -90 161 -86
rect 456 -88 460 -84
rect 466 -88 470 -84
rect 476 -88 480 -84
rect 486 -88 490 -84
rect 783 -85 787 -81
rect 793 -85 797 -81
rect 803 -85 807 -81
rect 813 -85 817 -81
rect 328 -204 332 -200
rect 358 -206 362 -202
rect 421 -204 425 -200
rect 451 -206 455 -202
rect 508 -204 512 -200
rect 339 -216 343 -212
rect 538 -206 542 -202
rect 432 -216 436 -212
rect 519 -216 523 -212
<< pdcontact >>
rect 113 167 117 171
rect 123 174 127 178
rect 123 167 127 171
rect 133 169 137 173
rect 143 181 147 185
rect 143 174 147 178
rect 200 167 204 171
rect 210 174 214 178
rect 210 167 214 171
rect 220 169 224 173
rect 230 181 234 185
rect 230 174 234 178
rect 293 167 297 171
rect 303 174 307 178
rect 303 167 307 171
rect 313 169 317 173
rect 323 181 327 185
rect 323 174 327 178
rect 533 183 537 187
rect 533 176 537 180
rect 626 183 630 187
rect 543 171 547 175
rect 553 176 557 180
rect 553 169 557 173
rect 626 176 630 180
rect 563 169 567 173
rect 713 183 717 187
rect 636 171 640 175
rect 646 176 650 180
rect 646 169 650 173
rect 713 176 717 180
rect 656 169 660 173
rect 723 171 727 175
rect 733 176 737 180
rect 733 169 737 173
rect 743 169 747 173
rect 35 113 39 117
rect 45 113 49 117
rect 55 113 59 117
rect 65 117 69 121
rect 121 114 125 118
rect 131 135 135 139
rect 131 128 135 132
rect 147 114 151 118
rect 157 121 161 125
rect 167 129 171 133
rect 205 114 209 118
rect 215 135 219 139
rect 215 128 219 132
rect 231 114 235 118
rect 241 121 245 125
rect 251 129 255 133
rect 267 113 271 117
rect 277 113 281 117
rect 287 113 291 117
rect 297 117 301 121
rect 364 115 368 119
rect 374 115 378 119
rect 384 115 388 119
rect 394 119 398 123
rect 450 116 454 120
rect 460 137 464 141
rect 460 130 464 134
rect 476 116 480 120
rect 486 123 490 127
rect 496 131 500 135
rect 534 116 538 120
rect 544 137 548 141
rect 544 130 548 134
rect 560 116 564 120
rect 570 123 574 127
rect 580 131 584 135
rect 596 115 600 119
rect 606 115 610 119
rect 616 115 620 119
rect 626 119 630 123
rect 691 118 695 122
rect 701 118 705 122
rect 711 118 715 122
rect 721 122 725 126
rect 777 119 781 123
rect 787 140 791 144
rect 787 133 791 137
rect 803 119 807 123
rect 813 126 817 130
rect 823 134 827 138
rect 861 119 865 123
rect 871 140 875 144
rect 871 133 875 137
rect 887 119 891 123
rect 897 126 901 130
rect 907 134 911 138
rect 923 118 927 122
rect 933 118 937 122
rect 943 118 947 122
rect 953 122 957 126
rect 128 18 132 22
rect 158 20 162 24
rect 457 20 461 24
rect 146 11 150 15
rect 487 22 491 26
rect 784 23 788 27
rect 475 13 479 17
rect 814 25 818 29
rect 802 16 806 20
rect 34 -33 38 -29
rect 44 -33 48 -29
rect 54 -33 58 -29
rect 64 -29 68 -25
rect 120 -32 124 -28
rect 130 -11 134 -7
rect 130 -18 134 -14
rect 146 -32 150 -28
rect 156 -25 160 -21
rect 166 -17 170 -13
rect 204 -32 208 -28
rect 214 -11 218 -7
rect 214 -18 218 -14
rect 230 -32 234 -28
rect 240 -25 244 -21
rect 250 -17 254 -13
rect 266 -33 270 -29
rect 276 -33 280 -29
rect 286 -33 290 -29
rect 296 -29 300 -25
rect 363 -31 367 -27
rect 373 -31 377 -27
rect 383 -31 387 -27
rect 393 -27 397 -23
rect 449 -30 453 -26
rect 459 -9 463 -5
rect 459 -16 463 -12
rect 475 -30 479 -26
rect 485 -23 489 -19
rect 495 -15 499 -11
rect 533 -30 537 -26
rect 543 -9 547 -5
rect 543 -16 547 -12
rect 559 -30 563 -26
rect 569 -23 573 -19
rect 579 -15 583 -11
rect 595 -31 599 -27
rect 605 -31 609 -27
rect 615 -31 619 -27
rect 625 -27 629 -23
rect 690 -28 694 -24
rect 700 -28 704 -24
rect 710 -28 714 -24
rect 720 -24 724 -20
rect 776 -27 780 -23
rect 786 -6 790 -2
rect 786 -13 790 -9
rect 802 -27 806 -23
rect 812 -20 816 -16
rect 822 -12 826 -8
rect 860 -27 864 -23
rect 870 -6 874 -2
rect 870 -13 874 -9
rect 886 -27 890 -23
rect 896 -20 900 -16
rect 906 -12 910 -8
rect 922 -28 926 -24
rect 932 -28 936 -24
rect 942 -28 946 -24
rect 952 -24 956 -20
rect 127 -128 131 -124
rect 157 -126 161 -122
rect 456 -126 460 -122
rect 145 -135 149 -131
rect 486 -124 490 -120
rect 783 -123 787 -119
rect 474 -133 478 -129
rect 813 -121 817 -117
rect 801 -130 805 -126
rect 328 -173 332 -169
rect 328 -180 332 -176
rect 338 -168 342 -164
rect 348 -166 352 -162
rect 348 -173 352 -169
rect 358 -166 362 -162
rect 421 -173 425 -169
rect 421 -180 425 -176
rect 431 -168 435 -164
rect 441 -166 445 -162
rect 441 -173 445 -169
rect 451 -166 455 -162
rect 508 -173 512 -169
rect 508 -180 512 -176
rect 518 -168 522 -164
rect 528 -166 532 -162
rect 528 -173 532 -169
rect 538 -166 542 -162
<< m2contact >>
rect 472 233 477 239
rect 108 224 113 229
rect 30 206 35 212
rect 108 200 112 204
rect 100 174 105 179
rect 196 200 200 204
rect 192 174 196 178
rect 289 200 293 204
rect 337 205 341 209
rect 513 205 518 210
rect 241 173 245 177
rect 285 174 289 178
rect 471 194 476 199
rect 567 202 571 206
rect 337 182 341 186
rect 514 182 519 187
rect 571 176 575 180
rect 337 165 341 169
rect 515 165 519 169
rect 602 175 606 180
rect 660 201 664 205
rect 747 201 751 205
rect 664 176 668 180
rect 677 178 681 182
rect 230 148 234 152
rect 267 149 272 153
rect 578 154 583 159
rect 613 154 617 159
rect 676 154 680 158
rect 690 153 694 157
rect 700 178 704 182
rect 752 176 757 180
rect 700 154 704 158
rect 58 128 62 132
rect 201 128 205 132
rect 34 100 38 104
rect 66 102 70 106
rect 103 102 107 106
rect 123 101 127 105
rect 170 101 174 105
rect 207 101 211 105
rect 290 128 294 132
rect 259 85 263 89
rect 298 103 302 107
rect 15 74 19 78
rect 300 75 306 81
rect 127 33 131 37
rect 118 25 122 29
rect 320 51 324 55
rect 387 130 391 134
rect 530 130 534 134
rect 363 102 367 106
rect 395 104 399 108
rect 432 104 436 108
rect 452 103 456 107
rect 587 123 591 127
rect 499 103 503 107
rect 536 103 540 107
rect 619 130 623 134
rect 588 87 592 91
rect 627 105 631 109
rect 340 74 347 81
rect 627 77 633 83
rect 345 51 349 55
rect 417 51 421 55
rect 456 35 460 39
rect 447 27 451 31
rect 639 48 643 52
rect 714 133 718 137
rect 857 133 861 137
rect 749 123 753 127
rect 690 105 694 109
rect 722 107 726 111
rect 759 107 763 111
rect 779 106 783 110
rect 834 125 838 129
rect 826 106 830 110
rect 750 90 754 94
rect 835 90 839 94
rect 912 126 917 130
rect 863 106 867 110
rect 946 133 950 137
rect 915 90 919 94
rect 954 108 958 112
rect 667 76 674 83
rect 751 60 756 65
rect 671 48 675 52
rect 742 48 746 52
rect 300 3 305 7
rect 320 2 325 7
rect 764 53 768 57
rect 783 38 787 42
rect 774 30 778 34
rect 827 53 831 57
rect 835 47 839 52
rect 764 22 768 26
rect 752 16 756 20
rect 834 12 839 19
rect 57 -18 61 -14
rect 33 -46 37 -42
rect 65 -44 69 -40
rect 102 -44 106 -40
rect 122 -45 126 -41
rect 169 -45 173 -41
rect 200 -18 204 -14
rect 206 -45 210 -41
rect 183 -61 187 -57
rect 289 -18 293 -14
rect 258 -61 262 -57
rect 297 -43 301 -39
rect 300 -71 308 -64
rect 249 -81 253 -77
rect 126 -113 130 -109
rect 117 -121 121 -117
rect 244 -100 250 -94
rect 273 -100 278 -95
rect 298 -100 303 -95
rect 319 -100 324 -95
rect 386 -16 390 -12
rect 529 -16 533 -12
rect 422 -35 426 -31
rect 362 -44 366 -40
rect 394 -42 398 -38
rect 431 -42 435 -38
rect 451 -43 455 -39
rect 498 -43 502 -39
rect 422 -59 426 -55
rect 535 -43 539 -39
rect 618 -16 622 -12
rect 587 -59 591 -55
rect 626 -41 630 -37
rect 337 -71 342 -66
rect 627 -70 631 -66
rect 422 -85 426 -81
rect 422 -103 426 -99
rect 455 -111 459 -107
rect 446 -119 450 -115
rect 512 -93 518 -88
rect 600 -93 605 -88
rect 713 -13 717 -9
rect 856 -13 860 -9
rect 689 -41 693 -37
rect 721 -39 725 -35
rect 758 -39 762 -35
rect 778 -40 782 -36
rect 825 -40 829 -36
rect 862 -40 866 -36
rect 945 -13 949 -9
rect 914 -56 918 -52
rect 953 -38 957 -34
rect 667 -70 671 -66
rect 725 -79 729 -75
rect 664 -93 669 -88
rect 698 -93 703 -88
rect 495 -126 500 -121
rect 394 -133 398 -129
rect 782 -108 786 -104
rect 773 -116 777 -112
rect 830 -91 836 -86
rect 725 -120 729 -116
rect 394 -162 398 -158
rect 366 -199 371 -194
rect 386 -210 390 -206
rect 496 -170 500 -165
rect 463 -182 467 -177
rect 459 -199 464 -194
rect 552 -182 556 -178
rect 544 -199 549 -194
rect 310 -221 317 -214
<< m3contact >>
rect 496 150 500 154
rect 515 129 519 133
<< psubstratepcontact >>
rect 142 217 146 221
rect 229 217 233 221
rect 322 217 326 221
rect 534 219 538 223
rect 627 219 631 223
rect 714 219 718 223
rect 36 78 40 82
rect 114 78 118 82
rect 198 78 202 82
rect 268 78 272 82
rect 365 80 369 84
rect 443 80 447 84
rect 527 80 531 84
rect 597 80 601 84
rect 692 83 696 87
rect 770 83 774 87
rect 854 83 858 87
rect 924 83 928 87
rect 129 68 133 72
rect 157 68 161 72
rect 458 70 462 74
rect 486 70 490 74
rect 785 73 789 77
rect 813 73 817 77
rect 35 -68 39 -64
rect 113 -68 117 -64
rect 197 -68 201 -64
rect 267 -68 271 -64
rect 364 -66 368 -62
rect 442 -66 446 -62
rect 526 -66 530 -62
rect 596 -66 600 -62
rect 691 -63 695 -59
rect 769 -63 773 -59
rect 853 -63 857 -59
rect 923 -63 927 -59
rect 128 -78 132 -74
rect 156 -78 160 -74
rect 457 -76 461 -72
rect 485 -76 489 -72
rect 784 -73 788 -69
rect 812 -73 816 -69
rect 329 -216 333 -212
rect 422 -216 426 -212
rect 509 -216 513 -212
<< nsubstratencontact >>
rect 142 157 146 161
rect 229 157 233 161
rect 322 157 326 161
rect 534 159 538 163
rect 627 159 631 163
rect 714 159 718 163
rect 36 138 40 142
rect 50 138 54 142
rect 64 138 68 142
rect 147 138 151 142
rect 231 138 235 142
rect 268 138 272 142
rect 282 138 286 142
rect 296 138 300 142
rect 365 140 369 144
rect 379 140 383 144
rect 393 140 397 144
rect 476 140 480 144
rect 560 140 564 144
rect 597 140 601 144
rect 611 140 615 144
rect 625 140 629 144
rect 692 143 696 147
rect 706 143 710 147
rect 720 143 724 147
rect 803 143 807 147
rect 887 143 891 147
rect 924 143 928 147
rect 938 143 942 147
rect 952 143 956 147
rect 157 8 161 12
rect 486 10 490 14
rect 813 13 817 17
rect 35 -8 39 -4
rect 49 -8 53 -4
rect 63 -8 67 -4
rect 146 -8 150 -4
rect 230 -8 234 -4
rect 267 -8 271 -4
rect 281 -8 285 -4
rect 295 -8 299 -4
rect 364 -6 368 -2
rect 378 -6 382 -2
rect 392 -6 396 -2
rect 475 -6 479 -2
rect 559 -6 563 -2
rect 596 -6 600 -2
rect 610 -6 614 -2
rect 624 -6 628 -2
rect 691 -3 695 1
rect 705 -3 709 1
rect 719 -3 723 1
rect 802 -3 806 1
rect 886 -3 890 1
rect 923 -3 927 1
rect 937 -3 941 1
rect 951 -3 955 1
rect 156 -138 160 -134
rect 485 -136 489 -132
rect 812 -133 816 -129
rect 329 -156 333 -152
rect 422 -156 426 -152
rect 509 -156 513 -152
<< psubstratepdiff >>
rect 533 223 539 224
rect 141 221 147 222
rect 141 217 142 221
rect 146 217 147 221
rect 141 216 147 217
rect 228 221 234 222
rect 228 217 229 221
rect 233 217 234 221
rect 228 216 234 217
rect 321 221 327 222
rect 321 217 322 221
rect 326 217 327 221
rect 533 219 534 223
rect 538 219 539 223
rect 533 218 539 219
rect 626 223 632 224
rect 626 219 627 223
rect 631 219 632 223
rect 321 216 327 217
rect 626 218 632 219
rect 713 223 719 224
rect 713 219 714 223
rect 718 219 719 223
rect 713 218 719 219
rect 35 82 41 83
rect 35 78 36 82
rect 40 78 41 82
rect 35 77 41 78
rect 113 82 119 83
rect 113 78 114 82
rect 118 78 119 82
rect 113 77 119 78
rect 197 82 203 83
rect 197 78 198 82
rect 202 78 203 82
rect 197 77 203 78
rect 364 84 370 85
rect 267 82 273 83
rect 267 78 268 82
rect 272 78 273 82
rect 267 77 273 78
rect 364 80 365 84
rect 369 80 370 84
rect 364 79 370 80
rect 442 84 448 85
rect 442 80 443 84
rect 447 80 448 84
rect 442 79 448 80
rect 526 84 532 85
rect 526 80 527 84
rect 531 80 532 84
rect 526 79 532 80
rect 691 87 697 88
rect 596 84 602 85
rect 596 80 597 84
rect 601 80 602 84
rect 596 79 602 80
rect 691 83 692 87
rect 696 83 697 87
rect 691 82 697 83
rect 769 87 775 88
rect 769 83 770 87
rect 774 83 775 87
rect 769 82 775 83
rect 853 87 859 88
rect 853 83 854 87
rect 858 83 859 87
rect 853 82 859 83
rect 923 87 929 88
rect 923 83 924 87
rect 928 83 929 87
rect 923 82 929 83
rect 784 77 818 78
rect 457 74 491 75
rect 128 72 162 73
rect 128 68 129 72
rect 133 68 157 72
rect 161 68 162 72
rect 457 70 458 74
rect 462 70 486 74
rect 490 70 491 74
rect 784 73 785 77
rect 789 73 813 77
rect 817 73 818 77
rect 784 72 818 73
rect 457 69 491 70
rect 128 67 162 68
rect 34 -64 40 -63
rect 34 -68 35 -64
rect 39 -68 40 -64
rect 34 -69 40 -68
rect 112 -64 118 -63
rect 112 -68 113 -64
rect 117 -68 118 -64
rect 112 -69 118 -68
rect 196 -64 202 -63
rect 196 -68 197 -64
rect 201 -68 202 -64
rect 196 -69 202 -68
rect 363 -62 369 -61
rect 266 -64 272 -63
rect 266 -68 267 -64
rect 271 -68 272 -64
rect 266 -69 272 -68
rect 363 -66 364 -62
rect 368 -66 369 -62
rect 363 -67 369 -66
rect 441 -62 447 -61
rect 441 -66 442 -62
rect 446 -66 447 -62
rect 441 -67 447 -66
rect 525 -62 531 -61
rect 525 -66 526 -62
rect 530 -66 531 -62
rect 525 -67 531 -66
rect 690 -59 696 -58
rect 595 -62 601 -61
rect 595 -66 596 -62
rect 600 -66 601 -62
rect 595 -67 601 -66
rect 690 -63 691 -59
rect 695 -63 696 -59
rect 690 -64 696 -63
rect 768 -59 774 -58
rect 768 -63 769 -59
rect 773 -63 774 -59
rect 768 -64 774 -63
rect 852 -59 858 -58
rect 852 -63 853 -59
rect 857 -63 858 -59
rect 852 -64 858 -63
rect 922 -59 928 -58
rect 922 -63 923 -59
rect 927 -63 928 -59
rect 922 -64 928 -63
rect 783 -69 817 -68
rect 456 -72 490 -71
rect 127 -74 161 -73
rect 127 -78 128 -74
rect 132 -78 156 -74
rect 160 -78 161 -74
rect 456 -76 457 -72
rect 461 -76 485 -72
rect 489 -76 490 -72
rect 783 -73 784 -69
rect 788 -73 812 -69
rect 816 -73 817 -69
rect 783 -74 817 -73
rect 456 -77 490 -76
rect 127 -79 161 -78
rect 328 -212 334 -211
rect 328 -216 329 -212
rect 333 -216 334 -212
rect 328 -217 334 -216
rect 421 -212 427 -211
rect 421 -216 422 -212
rect 426 -216 427 -212
rect 421 -217 427 -216
rect 508 -212 514 -211
rect 508 -216 509 -212
rect 513 -216 514 -212
rect 508 -217 514 -216
<< nsubstratendiff >>
rect 141 161 147 162
rect 228 161 234 162
rect 533 163 539 164
rect 626 163 632 164
rect 713 163 719 164
rect 321 161 327 162
rect 141 157 142 161
rect 146 157 147 161
rect 141 156 147 157
rect 228 157 229 161
rect 233 157 234 161
rect 228 156 234 157
rect 321 157 322 161
rect 326 157 327 161
rect 533 159 534 163
rect 538 159 539 163
rect 533 158 539 159
rect 626 159 627 163
rect 631 159 632 163
rect 626 158 632 159
rect 713 159 714 163
rect 718 159 719 163
rect 713 158 719 159
rect 321 156 327 157
rect 364 144 398 145
rect 35 142 69 143
rect 35 138 36 142
rect 40 138 50 142
rect 54 138 64 142
rect 68 138 69 142
rect 146 142 152 143
rect 35 137 69 138
rect 146 138 147 142
rect 151 138 152 142
rect 230 142 236 143
rect 146 137 152 138
rect 230 138 231 142
rect 235 138 236 142
rect 267 142 301 143
rect 230 137 236 138
rect 267 138 268 142
rect 272 138 282 142
rect 286 138 296 142
rect 300 138 301 142
rect 364 140 365 144
rect 369 140 379 144
rect 383 140 393 144
rect 397 140 398 144
rect 475 144 481 145
rect 364 139 398 140
rect 267 137 301 138
rect 475 140 476 144
rect 480 140 481 144
rect 559 144 565 145
rect 475 139 481 140
rect 559 140 560 144
rect 564 140 565 144
rect 596 144 630 145
rect 559 139 565 140
rect 596 140 597 144
rect 601 140 611 144
rect 615 140 625 144
rect 629 140 630 144
rect 691 143 692 147
rect 696 143 706 147
rect 710 143 720 147
rect 724 143 725 147
rect 802 147 808 148
rect 691 142 725 143
rect 596 139 630 140
rect 802 143 803 147
rect 807 143 808 147
rect 886 147 892 148
rect 802 142 808 143
rect 886 143 887 147
rect 891 143 892 147
rect 923 147 957 148
rect 886 142 892 143
rect 923 143 924 147
rect 928 143 938 147
rect 942 143 952 147
rect 956 143 957 147
rect 923 142 957 143
rect 156 12 162 13
rect 812 17 818 18
rect 485 14 491 15
rect 156 8 157 12
rect 161 8 162 12
rect 485 10 486 14
rect 490 10 491 14
rect 812 13 813 17
rect 817 13 818 17
rect 812 12 818 13
rect 485 9 491 10
rect 156 7 162 8
rect 690 1 724 2
rect 363 -2 397 -1
rect 34 -4 68 -3
rect 34 -8 35 -4
rect 39 -8 49 -4
rect 53 -8 63 -4
rect 67 -8 68 -4
rect 145 -4 151 -3
rect 34 -9 68 -8
rect 145 -8 146 -4
rect 150 -8 151 -4
rect 229 -4 235 -3
rect 145 -9 151 -8
rect 229 -8 230 -4
rect 234 -8 235 -4
rect 266 -4 300 -3
rect 229 -9 235 -8
rect 266 -8 267 -4
rect 271 -8 281 -4
rect 285 -8 295 -4
rect 299 -8 300 -4
rect 363 -6 364 -2
rect 368 -6 378 -2
rect 382 -6 392 -2
rect 396 -6 397 -2
rect 474 -2 480 -1
rect 363 -7 397 -6
rect 266 -9 300 -8
rect 474 -6 475 -2
rect 479 -6 480 -2
rect 558 -2 564 -1
rect 474 -7 480 -6
rect 558 -6 559 -2
rect 563 -6 564 -2
rect 595 -2 629 -1
rect 558 -7 564 -6
rect 595 -6 596 -2
rect 600 -6 610 -2
rect 614 -6 624 -2
rect 628 -6 629 -2
rect 690 -3 691 1
rect 695 -3 705 1
rect 709 -3 719 1
rect 723 -3 724 1
rect 801 1 807 2
rect 690 -4 724 -3
rect 595 -7 629 -6
rect 801 -3 802 1
rect 806 -3 807 1
rect 885 1 891 2
rect 801 -4 807 -3
rect 885 -3 886 1
rect 890 -3 891 1
rect 922 1 956 2
rect 885 -4 891 -3
rect 922 -3 923 1
rect 927 -3 937 1
rect 941 -3 951 1
rect 955 -3 956 1
rect 922 -4 956 -3
rect 155 -134 161 -133
rect 811 -129 817 -128
rect 484 -132 490 -131
rect 155 -138 156 -134
rect 160 -138 161 -134
rect 484 -136 485 -132
rect 489 -136 490 -132
rect 811 -133 812 -129
rect 816 -133 817 -129
rect 811 -134 817 -133
rect 484 -137 490 -136
rect 155 -139 161 -138
rect 328 -152 334 -151
rect 328 -156 329 -152
rect 333 -156 334 -152
rect 421 -152 427 -151
rect 421 -156 422 -152
rect 426 -156 427 -152
rect 508 -152 514 -151
rect 508 -156 509 -152
rect 513 -156 514 -152
rect 328 -157 334 -156
rect 421 -157 427 -156
rect 508 -157 514 -156
<< pad >>
rect 169 151 173 155
<< labels >>
rlabel metal1 474 74 474 74 2 vss
rlabel metal1 708 83 708 83 6 vss
rlabel metal1 940 147 940 147 6 vdd
rlabel metal1 801 77 801 77 2 vss
rlabel metal1 801 13 801 13 2 vdd
rlabel metal1 800 -133 800 -133 2 vdd
rlabel metal1 800 -69 800 -69 2 vss
rlabel metal1 939 -63 939 -63 6 vss
rlabel metal1 939 1 939 1 6 vdd
rlabel metal1 707 1 707 1 6 vdd
rlabel metal1 707 -63 707 -63 6 vss
rlabel metal1 797 1 797 1 6 vdd
rlabel metal1 473 -72 473 -72 2 vss
rlabel metal1 612 -66 612 -66 6 vss
rlabel metal1 612 -2 612 -2 6 vdd
rlabel metal1 380 -2 380 -2 6 vdd
rlabel metal1 380 -66 380 -66 6 vss
rlabel metal1 554 -2 554 -2 6 vdd
rlabel metal1 554 -66 554 -66 6 vss
rlabel metal1 144 -138 144 -138 2 vdd
rlabel metal1 51 -4 51 -4 6 vdd
rlabel metal1 51 -68 51 -68 6 vss
rlabel metal1 225 -4 225 -4 6 vdd
rlabel metal1 225 -68 225 -68 6 vss
rlabel m2contact 110 201 110 201 1 q0_M1
rlabel metal1 146 193 146 193 1 q0b2_M1
rlabel metal1 318 200 318 200 1 q0b0_n_M1
rlabel metal1 438 206 438 206 1 b2_M1
rlabel metal1 439 185 439 185 1 b1_M1
rlabel metal1 439 166 439 166 1 b0_M1
rlabel metal1 533 204 533 204 1 q1b0_M1
rlabel metal1 635 211 635 211 1 q1b1_M1
rlabel metal1 635 189 635 189 1 q1b1_n_M1
rlabel metal1 713 200 713 200 1 q1b2_M1
rlabel metal1 722 200 722 200 1 q1b2_n_M1
rlabel m2contact 749 203 749 203 1 q1_M1
rlabel metal1 938 111 938 111 1 zc1_n_3_M1
rlabel metal1 924 111 924 111 1 c1_3_M1
rlabel metal1 910 115 910 115 1 s_fa3_M1
rlabel metal1 887 133 887 133 1 cn_3_M1
rlabel ntransistor 903 98 903 98 1 s_fa3_n_M1
rlabel metal1 826 115 826 115 1 so_3_M1
rlabel metal1 814 136 814 136 1 bn3_M1
rlabel ptransistor 810 120 810 120 1 an3_M1
rlabel metal1 713 115 713 115 1 co_n3_M1
rlabel metal1 700 95 700 95 1 co_3_M1
rlabel metal1 597 108 597 108 1 c1_2_M1
rlabel metal1 611 108 611 108 1 zc1_2_n_M1
rlabel ntransistor 576 95 576 95 1 son_2_M1
rlabel pdcontact 573 125 573 125 1 s_fa2_M1
rlabel metal1 561 108 561 108 1 cn2_M1
rlabel metal1 499 112 499 112 1 so_2_M1
rlabel polycontact 489 108 489 108 1 an_2_M1
rlabel polycontact 483 109 483 109 1 bn_2_M1
rlabel metal1 386 111 386 111 1 co_n2_M1
rlabel metal1 373 92 373 92 1 co_2_M1
rlabel metal1 282 106 282 106 1 zc1_n1_M1
rlabel metal1 268 106 268 106 1 c1_1_M1
rlabel metal1 254 110 254 110 1 a1_M1
rlabel ntransistor 247 93 247 93 1 a1_n_M1
rlabel ntransistor 163 94 163 94 1 an_1_M1
rlabel metal1 170 110 170 110 1 so_1_M1
rlabel metal1 158 131 158 131 1 bn_1_M1
rlabel metal1 57 110 57 110 1 co_n1_M1
rlabel metal1 44 90 44 90 1 co_1_M1
rlabel metal1 153 38 153 38 1 c_fa1_n_M1
rlabel metal1 161 38 161 38 1 c_fa1_M1
rlabel metal1 482 42 482 42 1 c_fa_n_M1
rlabel metal1 490 46 490 46 1 c_fa2_M1
rlabel metal1 809 45 809 45 1 c_fa3_n_M1
rlabel metal1 817 49 817 49 1 c_fa3_M1
rlabel metal1 937 -35 937 -35 1 zc1_6_n_M1
rlabel metal1 923 -35 923 -35 1 c1_6_M1
rlabel ntransistor 902 -48 902 -48 1 s_fa_6_n_M1
rlabel metal1 909 -31 909 -31 1 a2_M1
rlabel metal1 885 -14 885 -14 1 cn_6_M1
rlabel metal1 825 -31 825 -31 1 so_6_M1
rlabel ptransistor 809 -26 809 -26 1 an_6_M1
rlabel metal1 770 -37 770 -37 1 bn_6_M1
rlabel metal1 712 -31 712 -31 1 co_n_6_M1
rlabel metal1 699 -51 699 -51 1 co_6_M1
rlabel metal1 610 -38 610 -38 1 zc1_n_5_M1
rlabel metal1 596 -38 596 -38 1 c1_5_M1
rlabel metal1 558 -18 558 -18 1 cn_5_M1
rlabel metal1 582 -34 582 -34 1 a3_M1
rlabel ntransistor 575 -51 575 -51 1 s_fa5_n_M1
rlabel metal1 486 -13 486 -13 1 bn_5_M1
rlabel ptransistor 482 -29 482 -29 1 an_5_M1
rlabel metal1 498 -34 498 -34 1 so_5_M1
rlabel metal1 385 -34 385 -34 1 co_5__M1
rlabel metal1 281 -40 281 -40 1 zc1_4_M1
rlabel metal1 267 -40 267 -40 1 c1_4_M1
rlabel metal1 253 -36 253 -36 1 a4_M1
rlabel ntransistor 246 -53 246 -53 1 s_fa4_n_M1
rlabel metal1 229 -20 229 -20 1 cn_1_M1
rlabel metal1 146 -21 146 -21 1 bn4_M1
rlabel ptransistor 153 -31 153 -31 1 an4_M1
rlabel metal1 169 -36 169 -36 1 so_4_M1
rlabel metal1 56 -36 56 -36 1 co_n4_M1
rlabel metal1 43 -56 43 -56 1 co_4_M1
rlabel metal1 152 -106 152 -106 1 a5_n_M1
rlabel metal1 160 -102 160 -102 1 a5_M1
rlabel metal1 489 -100 489 -100 1 c_fa5_M1
rlabel metal1 481 -104 481 -104 1 c_fa5_n_M1
rlabel metal1 808 -101 808 -101 1 c_fa6_n_M1
rlabel metal1 816 -97 816 -97 1 c_fa6_M1
rlabel metal1 509 -194 509 -194 1 q2b0_M1
rlabel metal1 518 -195 518 -195 1 q2b0_n_M1
rlabel m2contact 546 -196 546 -196 1 q2_M1
rlabel metal1 421 -194 421 -194 1 q2b1_M1
rlabel metal1 430 -194 430 -194 1 q2b1_n_M1
rlabel metal1 351 -205 351 -205 1 q2b2_n_M1
rlabel metal1 329 -206 329 -206 1 q2b2_M1
rlabel metal1 138 197 138 197 1 q0b2_n_M1
rlabel metal1 233 197 233 197 1 q0b1_M1
rlabel metal1 542 190 542 190 1 q1b0_n_M1
rlabel metal1 225 198 225 198 1 q0b1_n_M1
rlabel metal1 325 199 325 199 1 a0_M1
<< end >>
