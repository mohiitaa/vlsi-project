magic
tech scmos
timestamp 1523180881
<< pwell >>
rect 153 1041 171 1045
rect 151 1037 171 1041
rect 151 1001 199 1037
rect 238 1001 286 1037
rect 331 1001 379 1037
rect 571 1003 619 1039
rect 664 1003 712 1039
rect 751 1003 799 1039
rect 80 878 223 914
rect 235 878 353 914
rect 409 880 552 916
rect 564 880 682 916
rect 736 883 879 919
rect 1606 942 1642 1028
rect 891 883 1009 919
rect 166 852 214 878
rect 495 854 543 880
rect 822 857 870 883
rect 1580 894 1642 942
rect 1730 946 1766 1064
rect 1730 941 1754 946
rect 1732 934 1754 941
rect 1732 925 1766 934
rect 1606 885 1642 894
rect 1730 877 1792 925
rect 1413 829 1453 854
rect 1413 818 1454 829
rect 79 732 222 768
rect 234 732 352 768
rect 408 734 551 770
rect 563 734 681 770
rect 735 737 878 773
rect 1414 793 1454 818
rect 890 737 1008 773
rect 165 706 213 732
rect 494 708 542 734
rect 821 711 869 737
rect 1606 755 1642 873
rect 1730 791 1766 877
rect 2445 868 2493 894
rect 2672 870 2776 896
rect 2805 870 2853 896
rect 2306 832 2424 868
rect 1986 727 2129 752
rect 1413 678 1454 714
rect 1968 716 2129 727
rect 2436 832 2579 868
rect 2666 834 2784 870
rect 2796 834 2939 870
rect 2141 716 2259 752
rect 2342 742 2476 744
rect 2492 742 2615 744
rect 2342 720 2615 742
rect 366 584 414 620
rect 459 584 507 620
rect 546 584 594 620
rect 1608 582 1644 668
rect 164 535 182 539
rect 162 531 182 535
rect 1582 534 1644 582
rect 1732 586 1768 704
rect 1968 691 2120 716
rect 2342 708 2485 720
rect 2497 708 2615 720
rect 2702 744 2836 746
rect 2852 744 2975 746
rect 2702 722 2975 744
rect 2702 710 2845 722
rect 2857 710 2975 722
rect 2072 690 2120 691
rect 2428 682 2476 708
rect 2788 684 2836 710
rect 1732 581 1756 586
rect 1734 574 1756 581
rect 1734 565 1768 574
rect 162 495 210 531
rect 249 495 297 531
rect 342 495 390 531
rect 582 497 630 533
rect 675 497 723 533
rect 762 497 810 533
rect 1608 525 1644 534
rect 1732 517 1794 565
rect 91 372 234 408
rect 246 372 364 408
rect 420 374 563 410
rect 575 374 693 410
rect 747 377 890 413
rect 902 377 1020 413
rect 1608 395 1644 513
rect 1732 431 1768 517
rect 2029 464 2047 468
rect 2027 460 2047 464
rect 2027 424 2075 460
rect 2114 424 2162 460
rect 2207 424 2255 460
rect 2447 426 2495 462
rect 2540 426 2588 462
rect 2627 426 2675 462
rect 177 346 225 372
rect 506 348 554 374
rect 833 351 881 377
rect 1445 320 1485 356
rect 90 226 233 262
rect 245 226 363 262
rect 419 228 562 264
rect 574 228 692 264
rect 746 231 889 267
rect 901 231 1019 267
rect 176 200 224 226
rect 505 202 553 228
rect 832 205 880 231
rect 1724 230 1760 348
rect 1956 301 2099 337
rect 2111 301 2229 337
rect 2285 303 2428 339
rect 2440 303 2558 339
rect 2612 306 2755 342
rect 2767 306 2885 342
rect 2042 275 2090 301
rect 2371 277 2419 303
rect 2698 280 2746 306
rect 1447 187 1487 219
rect 1447 177 1488 187
rect 1447 175 1489 177
rect 377 78 425 114
rect 470 78 518 114
rect 1449 141 1489 175
rect 557 78 605 114
rect 1724 209 1760 218
rect 1724 166 1786 209
rect 1724 75 1785 166
rect 1749 57 1785 75
rect 1955 155 2098 191
rect 2110 155 2228 191
rect 2284 157 2427 193
rect 2439 157 2557 193
rect 2611 160 2754 196
rect 2766 160 2884 196
rect 2041 129 2089 155
rect 2370 131 2418 157
rect 2697 134 2745 160
rect 2242 7 2290 43
rect 2335 7 2383 43
rect 2422 7 2470 43
<< nwell >>
rect 1686 1063 1730 1064
rect 151 958 199 1001
rect 238 958 286 1001
rect 331 958 379 1001
rect 571 966 619 1003
rect 664 966 712 1003
rect 571 963 712 966
rect 567 960 712 963
rect 1048 1005 1227 1031
rect 1240 1005 1281 1031
rect 1296 1005 1337 1031
rect 1350 1005 1391 1031
rect 1679 1028 1730 1063
rect 751 972 799 1003
rect 751 963 812 972
rect 751 960 879 963
rect 80 914 223 958
rect 235 957 379 958
rect 235 914 353 957
rect 409 916 552 960
rect 564 946 879 960
rect 564 916 682 946
rect 736 919 879 946
rect 891 919 1009 963
rect 1560 942 1573 946
rect 1144 900 1231 926
rect 1244 900 1285 926
rect 1300 900 1341 926
rect 1354 900 1395 926
rect 166 845 214 852
rect 495 847 543 854
rect 1048 860 1227 886
rect 1240 860 1281 886
rect 1296 860 1337 886
rect 1350 860 1391 886
rect 822 850 870 857
rect 162 832 214 845
rect 491 834 543 847
rect 818 837 870 850
rect 166 816 214 832
rect 495 818 543 834
rect 822 824 870 837
rect 1413 854 1453 898
rect 1537 894 1580 942
rect 1642 941 1730 1028
rect 1642 925 1732 941
rect 1642 885 1730 925
rect 1682 873 1730 885
rect 1792 877 1836 925
rect 2445 914 2493 937
rect 2445 901 2497 914
rect 2445 894 2493 901
rect 155 812 221 816
rect 485 814 551 818
rect 793 817 904 824
rect 79 768 222 812
rect 234 768 352 812
rect 408 770 551 814
rect 563 770 681 814
rect 735 808 1008 817
rect 735 773 878 808
rect 890 773 1008 808
rect 1144 755 1231 781
rect 1244 755 1285 781
rect 1300 755 1341 781
rect 1354 758 1395 781
rect 1414 758 1454 793
rect 1383 755 1395 758
rect 165 699 213 706
rect 494 701 542 708
rect 1047 718 1226 744
rect 1239 718 1280 744
rect 1295 718 1336 744
rect 1349 718 1390 744
rect 821 704 869 711
rect 161 686 213 699
rect 490 688 542 701
rect 817 691 869 704
rect 165 662 213 686
rect 494 678 542 688
rect 368 664 600 678
rect 821 667 869 691
rect 1413 714 1454 758
rect 1642 791 1730 873
rect 1799 873 1812 877
rect 2672 896 2776 940
rect 2805 916 2853 939
rect 2805 903 2857 916
rect 2805 896 2853 903
rect 1642 757 1691 791
rect 1642 755 1686 757
rect 1986 752 2129 796
rect 2141 752 2259 796
rect 2306 792 2424 832
rect 2436 795 2579 832
rect 2436 792 2614 795
rect 2306 788 2614 792
rect 2666 794 2784 834
rect 2796 797 2939 834
rect 2796 794 2974 797
rect 2666 790 2974 794
rect 2308 783 2615 788
rect 2668 785 2975 790
rect 2342 744 2615 783
rect 2476 742 2492 744
rect 1688 703 1732 704
rect 1681 668 1732 703
rect 366 661 600 664
rect 366 620 414 661
rect 459 620 507 661
rect 546 620 594 661
rect 1143 613 1230 639
rect 1243 613 1284 639
rect 1299 613 1340 639
rect 1353 613 1394 639
rect 1562 582 1575 586
rect 1539 534 1582 582
rect 1644 581 1732 668
rect 2702 746 2975 785
rect 2836 744 2852 746
rect 1968 690 2072 691
rect 1968 647 2120 690
rect 2428 675 2476 682
rect 2788 677 2836 684
rect 2424 662 2476 675
rect 2784 664 2836 677
rect 2072 646 2120 647
rect 2428 638 2476 662
rect 2788 640 2836 664
rect 1644 565 1734 581
rect 162 452 210 495
rect 249 452 297 495
rect 342 452 390 495
rect 582 460 630 497
rect 675 460 723 497
rect 582 457 723 460
rect 578 454 723 457
rect 1644 525 1732 565
rect 762 466 810 497
rect 1069 494 1248 520
rect 1261 494 1302 520
rect 1317 494 1358 520
rect 1371 494 1412 520
rect 1684 513 1732 525
rect 1794 517 1838 565
rect 762 457 823 466
rect 762 454 890 457
rect 91 408 234 452
rect 246 451 390 452
rect 246 408 364 451
rect 420 410 563 454
rect 575 440 890 454
rect 575 410 693 440
rect 747 413 890 440
rect 902 413 1020 457
rect 1165 389 1252 415
rect 1265 389 1306 415
rect 1321 389 1362 415
rect 1375 389 1416 415
rect 1644 431 1732 513
rect 1801 513 1814 517
rect 1644 397 1693 431
rect 1644 395 1688 397
rect 2027 381 2075 424
rect 2114 381 2162 424
rect 2207 381 2255 424
rect 2447 389 2495 426
rect 2540 389 2588 426
rect 2447 386 2588 389
rect 2443 383 2588 386
rect 2627 395 2675 426
rect 2627 386 2688 395
rect 2627 383 2755 386
rect 177 339 225 346
rect 506 341 554 348
rect 833 344 881 351
rect 1067 349 1246 375
rect 1259 349 1300 375
rect 1315 349 1356 375
rect 1369 349 1410 375
rect 173 326 225 339
rect 502 328 554 341
rect 829 331 881 344
rect 177 310 225 326
rect 506 312 554 328
rect 833 318 881 331
rect 166 306 232 310
rect 496 308 562 312
rect 804 311 915 318
rect 90 262 233 306
rect 245 262 363 306
rect 419 264 562 308
rect 574 264 692 308
rect 746 302 1019 311
rect 746 267 889 302
rect 901 267 1019 302
rect 1445 279 1485 320
rect 1444 276 1485 279
rect 1163 244 1250 270
rect 1263 244 1304 270
rect 1319 244 1360 270
rect 1373 244 1414 270
rect 1444 263 1484 276
rect 176 193 224 200
rect 505 195 553 202
rect 1068 207 1247 233
rect 1260 207 1301 233
rect 1316 207 1357 233
rect 1370 207 1411 233
rect 1447 219 1487 263
rect 1680 230 1724 348
rect 1956 337 2099 381
rect 2111 380 2255 381
rect 2111 337 2229 380
rect 2285 339 2428 383
rect 2440 369 2755 383
rect 2440 339 2558 369
rect 2612 342 2755 369
rect 2767 342 2885 386
rect 2042 268 2090 275
rect 2371 270 2419 277
rect 2698 273 2746 280
rect 2038 255 2090 268
rect 2367 257 2419 270
rect 2694 260 2746 273
rect 2042 239 2090 255
rect 2371 241 2419 257
rect 2698 247 2746 260
rect 2031 235 2097 239
rect 2361 237 2427 241
rect 2669 240 2780 247
rect 832 198 880 205
rect 172 180 224 193
rect 501 182 553 195
rect 828 185 880 198
rect 176 156 224 180
rect 505 172 553 182
rect 379 158 611 172
rect 832 161 880 185
rect 377 155 611 158
rect 377 114 425 155
rect 470 114 518 155
rect 557 114 605 155
rect 1164 102 1251 128
rect 1264 102 1305 128
rect 1320 102 1361 128
rect 1374 102 1415 128
rect 1449 97 1489 141
rect 1680 75 1724 218
rect 1786 166 1830 209
rect 1785 161 1830 166
rect 1955 191 2098 235
rect 1785 57 1829 161
rect 2110 191 2228 235
rect 2284 193 2427 237
rect 2439 193 2557 237
rect 2611 231 2884 240
rect 2611 196 2754 231
rect 2766 196 2884 231
rect 2041 122 2089 129
rect 2370 124 2418 131
rect 2697 127 2745 134
rect 2037 109 2089 122
rect 2366 111 2418 124
rect 2693 114 2745 127
rect 2041 85 2089 109
rect 2370 101 2418 111
rect 2244 87 2476 101
rect 2697 90 2745 114
rect 2242 84 2476 87
rect 2242 43 2290 84
rect 2335 43 2383 84
rect 2422 43 2470 84
<< polysilicon >>
rect 1735 1053 1741 1054
rect 1735 1051 1736 1053
rect 1709 1049 1714 1051
rect 1724 1049 1736 1051
rect 1740 1050 1741 1053
rect 1740 1049 1744 1050
rect 1735 1048 1744 1049
rect 1753 1048 1758 1050
rect 1703 1044 1709 1045
rect 1703 1040 1704 1044
rect 1708 1041 1709 1044
rect 1727 1041 1744 1043
rect 1753 1041 1758 1043
rect 1708 1040 1714 1041
rect 1703 1039 1714 1040
rect 1724 1039 1730 1041
rect 164 1020 166 1025
rect 171 1020 173 1025
rect 184 1018 186 1022
rect 251 1020 253 1025
rect 258 1020 260 1025
rect 271 1018 273 1022
rect 344 1020 346 1025
rect 351 1020 353 1025
rect 364 1018 366 1022
rect 584 1020 586 1024
rect 597 1022 599 1027
rect 604 1022 606 1027
rect 677 1020 679 1024
rect 690 1022 692 1027
rect 697 1022 699 1027
rect 764 1020 766 1024
rect 777 1022 779 1027
rect 784 1022 786 1027
rect 1085 1018 1087 1020
rect 1157 1018 1159 1024
rect 1196 1018 1198 1024
rect 1217 1018 1219 1024
rect 1250 1018 1252 1024
rect 1271 1018 1273 1024
rect 1306 1018 1308 1024
rect 1327 1018 1329 1024
rect 1360 1018 1362 1024
rect 1381 1018 1383 1024
rect 1727 1034 1733 1035
rect 1727 1031 1728 1034
rect 1707 1029 1712 1031
rect 1724 1030 1728 1031
rect 1732 1031 1733 1034
rect 1732 1030 1741 1031
rect 1724 1029 1741 1030
rect 1747 1029 1751 1031
rect 1621 1020 1625 1022
rect 1631 1021 1648 1022
rect 1631 1020 1640 1021
rect 1639 1017 1640 1020
rect 1644 1020 1648 1021
rect 1660 1020 1665 1022
rect 1644 1017 1645 1020
rect 1639 1016 1645 1017
rect 164 996 166 1009
rect 171 1004 173 1009
rect 184 1004 186 1009
rect 170 1003 176 1004
rect 170 999 171 1003
rect 175 999 176 1003
rect 170 998 176 999
rect 180 1003 186 1004
rect 180 999 181 1003
rect 185 999 186 1003
rect 180 998 186 999
rect 160 995 166 996
rect 160 991 161 995
rect 165 991 166 995
rect 160 990 166 991
rect 164 987 166 990
rect 174 987 176 998
rect 184 994 186 998
rect 251 996 253 1009
rect 258 1004 260 1009
rect 271 1004 273 1009
rect 257 1003 263 1004
rect 257 999 258 1003
rect 262 999 263 1003
rect 257 998 263 999
rect 267 1003 273 1004
rect 267 999 268 1003
rect 272 999 273 1003
rect 267 998 273 999
rect 247 995 253 996
rect 247 991 248 995
rect 252 991 253 995
rect 247 990 253 991
rect 251 987 253 990
rect 261 987 263 998
rect 271 994 273 998
rect 344 996 346 1009
rect 351 1004 353 1009
rect 364 1004 366 1009
rect 350 1003 356 1004
rect 350 999 351 1003
rect 355 999 356 1003
rect 350 998 356 999
rect 360 1003 366 1004
rect 360 999 361 1003
rect 365 999 366 1003
rect 360 998 366 999
rect 340 995 346 996
rect 164 969 166 974
rect 174 969 176 974
rect 184 972 186 976
rect 340 991 341 995
rect 345 991 346 995
rect 340 990 346 991
rect 344 987 346 990
rect 354 987 356 998
rect 364 994 366 998
rect 584 1006 586 1011
rect 597 1006 599 1011
rect 584 1005 590 1006
rect 584 1001 585 1005
rect 589 1001 590 1005
rect 584 1000 590 1001
rect 594 1005 600 1006
rect 594 1001 595 1005
rect 599 1001 600 1005
rect 594 1000 600 1001
rect 584 996 586 1000
rect 251 969 253 974
rect 261 969 263 974
rect 271 972 273 976
rect 594 989 596 1000
rect 604 998 606 1011
rect 677 1006 679 1011
rect 690 1006 692 1011
rect 677 1005 683 1006
rect 677 1001 678 1005
rect 682 1001 683 1005
rect 677 1000 683 1001
rect 687 1005 693 1006
rect 687 1001 688 1005
rect 692 1001 693 1005
rect 687 1000 693 1001
rect 604 997 610 998
rect 604 993 605 997
rect 609 993 610 997
rect 677 996 679 1000
rect 604 992 610 993
rect 604 989 606 992
rect 344 969 346 974
rect 354 969 356 974
rect 364 972 366 976
rect 584 974 586 978
rect 687 989 689 1000
rect 697 998 699 1011
rect 764 1006 766 1011
rect 777 1006 779 1011
rect 764 1005 770 1006
rect 764 1001 765 1005
rect 769 1001 770 1005
rect 764 1000 770 1001
rect 774 1005 780 1006
rect 774 1001 775 1005
rect 779 1001 780 1005
rect 774 1000 780 1001
rect 697 997 703 998
rect 697 993 698 997
rect 702 993 703 997
rect 764 996 766 1000
rect 697 992 703 993
rect 697 989 699 992
rect 594 971 596 976
rect 604 971 606 976
rect 677 974 679 978
rect 774 989 776 1000
rect 784 998 786 1011
rect 1085 1001 1087 1012
rect 784 997 790 998
rect 1157 1000 1159 1012
rect 1196 1000 1198 1012
rect 1217 1000 1219 1012
rect 1250 1000 1252 1012
rect 1271 1000 1273 1012
rect 1306 1000 1308 1012
rect 1327 1000 1329 1012
rect 1360 1000 1362 1012
rect 1381 1000 1383 1012
rect 1642 1010 1648 1012
rect 1658 1011 1669 1012
rect 1658 1010 1664 1011
rect 1614 1008 1619 1010
rect 1628 1008 1645 1010
rect 1663 1007 1664 1010
rect 1668 1007 1669 1011
rect 1663 1006 1669 1007
rect 1614 1001 1619 1003
rect 1628 1002 1637 1003
rect 1628 1001 1632 1002
rect 784 993 785 997
rect 789 993 790 997
rect 784 992 790 993
rect 784 989 786 992
rect 687 971 689 976
rect 697 971 699 976
rect 764 974 766 978
rect 1085 979 1087 997
rect 1197 996 1198 1000
rect 1218 996 1219 1000
rect 1251 996 1252 1000
rect 1272 996 1273 1000
rect 1307 996 1308 1000
rect 1328 996 1329 1000
rect 1361 996 1362 1000
rect 1382 996 1383 1000
rect 774 971 776 976
rect 784 971 786 976
rect 1085 973 1087 976
rect 1157 978 1159 996
rect 1196 981 1198 996
rect 1217 981 1219 996
rect 1250 981 1252 996
rect 1271 981 1273 996
rect 1306 981 1308 996
rect 1327 981 1329 996
rect 1360 981 1362 996
rect 1381 981 1383 996
rect 1631 998 1632 1001
rect 1636 1000 1648 1002
rect 1658 1000 1663 1002
rect 1636 998 1637 1000
rect 1631 997 1637 998
rect 1692 1003 1696 1005
rect 1723 1004 1732 1005
rect 1723 1003 1727 1004
rect 1726 1000 1727 1003
rect 1731 1002 1741 1004
rect 1753 1002 1758 1004
rect 1731 1000 1732 1002
rect 1726 999 1732 1000
rect 1736 995 1741 997
rect 1753 995 1758 997
rect 1701 993 1705 995
rect 1723 994 1738 995
rect 1723 993 1727 994
rect 1726 990 1727 993
rect 1731 993 1738 994
rect 1731 990 1732 993
rect 1726 989 1732 990
rect 1736 985 1741 987
rect 1750 985 1760 987
rect 1701 983 1705 985
rect 1723 983 1728 985
rect 1726 977 1728 983
rect 1726 975 1741 977
rect 1750 975 1754 977
rect 1157 972 1159 975
rect 1196 972 1198 975
rect 1217 972 1219 975
rect 1250 972 1252 975
rect 1271 972 1273 975
rect 1306 972 1308 975
rect 1327 972 1329 975
rect 1360 972 1362 975
rect 1381 972 1383 975
rect 1732 973 1738 975
rect 1732 969 1733 973
rect 1737 969 1738 973
rect 1692 967 1696 969
rect 1723 967 1728 969
rect 1732 968 1738 969
rect 1726 961 1728 967
rect 1758 964 1760 985
rect 1748 962 1760 964
rect 1748 961 1750 962
rect 1726 959 1736 961
rect 1745 959 1750 961
rect 172 948 174 952
rect 96 940 102 941
rect 86 932 88 937
rect 96 936 97 940
rect 101 936 102 940
rect 96 935 102 936
rect 96 930 98 935
rect 106 930 108 935
rect 157 932 163 933
rect 157 928 158 932
rect 162 928 163 932
rect 157 927 163 928
rect 86 917 88 920
rect 96 917 98 920
rect 86 916 92 917
rect 86 912 87 916
rect 91 912 92 916
rect 96 914 100 917
rect 86 911 92 912
rect 86 903 88 911
rect 98 900 100 914
rect 106 909 108 920
rect 161 918 163 927
rect 208 948 210 952
rect 256 948 258 952
rect 188 939 190 943
rect 198 939 200 943
rect 241 932 247 933
rect 241 928 242 932
rect 246 928 247 932
rect 241 927 247 928
rect 172 918 174 921
rect 188 918 190 921
rect 198 918 200 921
rect 208 918 210 921
rect 161 916 174 918
rect 180 916 190 918
rect 194 917 200 918
rect 105 908 111 909
rect 164 908 166 916
rect 180 912 182 916
rect 194 913 195 917
rect 199 913 200 917
rect 194 912 200 913
rect 204 917 210 918
rect 204 913 205 917
rect 209 913 210 917
rect 245 918 247 927
rect 292 948 294 952
rect 272 939 274 943
rect 282 939 284 943
rect 501 950 503 954
rect 425 942 431 943
rect 328 940 334 941
rect 318 932 320 937
rect 328 936 329 940
rect 333 936 334 940
rect 328 935 334 936
rect 256 918 258 921
rect 272 918 274 921
rect 282 918 284 921
rect 292 918 294 921
rect 328 930 330 935
rect 338 930 340 935
rect 415 934 417 939
rect 425 938 426 942
rect 430 938 431 942
rect 425 937 431 938
rect 425 932 427 937
rect 435 932 437 937
rect 486 934 492 935
rect 486 930 487 934
rect 491 930 492 934
rect 486 929 492 930
rect 245 916 258 918
rect 264 916 274 918
rect 278 917 284 918
rect 204 912 210 913
rect 173 911 182 912
rect 105 904 106 908
rect 110 904 111 908
rect 105 903 111 904
rect 105 900 107 903
rect 86 893 88 897
rect 173 907 174 911
rect 178 907 182 911
rect 198 908 200 912
rect 173 906 182 907
rect 180 903 182 906
rect 190 903 192 908
rect 198 906 202 908
rect 200 903 202 906
rect 207 903 209 912
rect 248 908 250 916
rect 264 912 266 916
rect 278 913 279 917
rect 283 913 284 917
rect 278 912 284 913
rect 288 917 294 918
rect 288 913 289 917
rect 293 913 294 917
rect 288 912 294 913
rect 318 917 320 920
rect 328 917 330 920
rect 318 916 324 917
rect 318 912 319 916
rect 323 912 324 916
rect 328 914 332 917
rect 257 911 266 912
rect 164 896 166 899
rect 164 894 169 896
rect 98 886 100 891
rect 105 886 107 891
rect 167 886 169 894
rect 180 890 182 894
rect 190 886 192 894
rect 257 907 258 911
rect 262 907 266 911
rect 282 908 284 912
rect 257 906 266 907
rect 264 903 266 906
rect 274 903 276 908
rect 282 906 286 908
rect 284 903 286 906
rect 291 903 293 912
rect 318 911 324 912
rect 318 903 320 911
rect 248 896 250 899
rect 248 894 253 896
rect 200 886 202 891
rect 207 886 209 891
rect 167 884 192 886
rect 251 886 253 894
rect 264 890 266 894
rect 274 886 276 894
rect 330 900 332 914
rect 338 909 340 920
rect 415 919 417 922
rect 425 919 427 922
rect 415 918 421 919
rect 415 914 416 918
rect 420 914 421 918
rect 425 916 429 919
rect 415 913 421 914
rect 337 908 343 909
rect 337 904 338 908
rect 342 904 343 908
rect 415 905 417 913
rect 337 903 343 904
rect 337 900 339 903
rect 318 893 320 897
rect 427 902 429 916
rect 435 911 437 922
rect 490 920 492 929
rect 537 950 539 954
rect 585 950 587 954
rect 517 941 519 945
rect 527 941 529 945
rect 570 934 576 935
rect 570 930 571 934
rect 575 930 576 934
rect 570 929 576 930
rect 501 920 503 923
rect 517 920 519 923
rect 527 920 529 923
rect 537 920 539 923
rect 490 918 503 920
rect 509 918 519 920
rect 523 919 529 920
rect 434 910 440 911
rect 493 910 495 918
rect 509 914 511 918
rect 523 915 524 919
rect 528 915 529 919
rect 523 914 529 915
rect 533 919 539 920
rect 533 915 534 919
rect 538 915 539 919
rect 574 920 576 929
rect 621 950 623 954
rect 601 941 603 945
rect 611 941 613 945
rect 828 953 830 957
rect 752 945 758 946
rect 657 942 663 943
rect 647 934 649 939
rect 657 938 658 942
rect 662 938 663 942
rect 657 937 663 938
rect 742 937 744 942
rect 752 941 753 945
rect 757 941 758 945
rect 752 940 758 941
rect 585 920 587 923
rect 601 920 603 923
rect 611 920 613 923
rect 621 920 623 923
rect 657 932 659 937
rect 667 932 669 937
rect 752 935 754 940
rect 762 935 764 940
rect 813 937 819 938
rect 813 933 814 937
rect 818 933 819 937
rect 813 932 819 933
rect 742 922 744 925
rect 752 922 754 925
rect 574 918 587 920
rect 593 918 603 920
rect 607 919 613 920
rect 533 914 539 915
rect 502 913 511 914
rect 434 906 435 910
rect 439 906 440 910
rect 434 905 440 906
rect 434 902 436 905
rect 415 895 417 899
rect 502 909 503 913
rect 507 909 511 913
rect 527 910 529 914
rect 502 908 511 909
rect 509 905 511 908
rect 519 905 521 910
rect 527 908 531 910
rect 529 905 531 908
rect 536 905 538 914
rect 577 910 579 918
rect 593 914 595 918
rect 607 915 608 919
rect 612 915 613 919
rect 607 914 613 915
rect 617 919 623 920
rect 617 915 618 919
rect 622 915 623 919
rect 617 914 623 915
rect 647 919 649 922
rect 657 919 659 922
rect 647 918 653 919
rect 647 914 648 918
rect 652 914 653 918
rect 657 916 661 919
rect 586 913 595 914
rect 493 898 495 901
rect 493 896 498 898
rect 284 886 286 891
rect 291 886 293 891
rect 251 884 276 886
rect 330 886 332 891
rect 337 886 339 891
rect 427 888 429 893
rect 434 888 436 893
rect 496 888 498 896
rect 509 892 511 896
rect 519 888 521 896
rect 586 909 587 913
rect 591 909 595 913
rect 611 910 613 914
rect 586 908 595 909
rect 593 905 595 908
rect 603 905 605 910
rect 611 908 615 910
rect 613 905 615 908
rect 620 905 622 914
rect 647 913 653 914
rect 647 905 649 913
rect 577 898 579 901
rect 577 896 582 898
rect 529 888 531 893
rect 536 888 538 893
rect 496 886 521 888
rect 580 888 582 896
rect 593 892 595 896
rect 603 888 605 896
rect 659 902 661 916
rect 667 911 669 922
rect 742 921 748 922
rect 742 917 743 921
rect 747 917 748 921
rect 752 919 756 922
rect 742 916 748 917
rect 666 910 672 911
rect 666 906 667 910
rect 671 906 672 910
rect 742 908 744 916
rect 666 905 672 906
rect 666 902 668 905
rect 754 905 756 919
rect 762 914 764 925
rect 817 923 819 932
rect 864 953 866 957
rect 912 953 914 957
rect 844 944 846 948
rect 854 944 856 948
rect 897 937 903 938
rect 897 933 898 937
rect 902 933 903 937
rect 897 932 903 933
rect 828 923 830 926
rect 844 923 846 926
rect 854 923 856 926
rect 864 923 866 926
rect 817 921 830 923
rect 836 921 846 923
rect 850 922 856 923
rect 761 913 767 914
rect 820 913 822 921
rect 836 917 838 921
rect 850 918 851 922
rect 855 918 856 922
rect 850 917 856 918
rect 860 922 866 923
rect 860 918 861 922
rect 865 918 866 922
rect 901 923 903 932
rect 948 953 950 957
rect 1161 956 1163 959
rect 1200 956 1202 959
rect 1221 956 1223 959
rect 1254 956 1256 959
rect 1275 956 1277 959
rect 1310 956 1312 959
rect 1331 956 1333 959
rect 1364 956 1366 959
rect 1385 956 1387 959
rect 1726 958 1728 959
rect 1711 957 1728 958
rect 928 944 930 948
rect 938 944 940 948
rect 984 945 990 946
rect 974 937 976 942
rect 984 941 985 945
rect 989 941 990 945
rect 984 940 990 941
rect 912 923 914 926
rect 928 923 930 926
rect 938 923 940 926
rect 948 923 950 926
rect 984 935 986 940
rect 994 935 996 940
rect 1161 935 1163 953
rect 1711 953 1712 957
rect 1716 956 1728 957
rect 1716 953 1717 956
rect 1711 952 1717 953
rect 1200 935 1202 950
rect 1221 935 1223 950
rect 1254 935 1256 950
rect 1275 935 1277 950
rect 1310 935 1312 950
rect 1331 935 1333 950
rect 1364 935 1366 950
rect 1385 935 1387 950
rect 1655 950 1661 951
rect 1655 947 1656 950
rect 1644 946 1656 947
rect 1660 946 1661 950
rect 1644 945 1661 946
rect 1644 944 1646 945
rect 1622 942 1627 944
rect 1636 942 1646 944
rect 1622 941 1624 942
rect 1612 939 1624 941
rect 1201 931 1202 935
rect 1222 931 1223 935
rect 1255 931 1256 935
rect 1276 931 1277 935
rect 1311 931 1312 935
rect 1332 931 1333 935
rect 1365 931 1366 935
rect 1386 931 1387 935
rect 901 921 914 923
rect 920 921 930 923
rect 934 922 940 923
rect 860 917 866 918
rect 829 916 838 917
rect 761 909 762 913
rect 766 909 767 913
rect 761 908 767 909
rect 761 905 763 908
rect 647 895 649 899
rect 742 898 744 902
rect 829 912 830 916
rect 834 912 838 916
rect 854 913 856 917
rect 829 911 838 912
rect 836 908 838 911
rect 846 908 848 913
rect 854 911 858 913
rect 856 908 858 911
rect 863 908 865 917
rect 904 913 906 921
rect 920 917 922 921
rect 934 918 935 922
rect 939 918 940 922
rect 934 917 940 918
rect 944 922 950 923
rect 944 918 945 922
rect 949 918 950 922
rect 944 917 950 918
rect 974 922 976 925
rect 984 922 986 925
rect 974 921 980 922
rect 974 917 975 921
rect 979 917 980 921
rect 984 919 988 922
rect 913 916 922 917
rect 820 901 822 904
rect 820 899 825 901
rect 613 888 615 893
rect 620 888 622 893
rect 580 886 605 888
rect 659 888 661 893
rect 666 888 668 893
rect 754 891 756 896
rect 761 891 763 896
rect 823 891 825 899
rect 836 895 838 899
rect 846 891 848 899
rect 913 912 914 916
rect 918 912 922 916
rect 938 913 940 917
rect 913 911 922 912
rect 920 908 922 911
rect 930 908 932 913
rect 938 911 942 913
rect 940 908 942 911
rect 947 908 949 917
rect 974 916 980 917
rect 974 908 976 916
rect 904 901 906 904
rect 904 899 909 901
rect 856 891 858 896
rect 863 891 865 896
rect 823 889 848 891
rect 907 891 909 899
rect 920 895 922 899
rect 930 891 932 899
rect 986 905 988 919
rect 994 914 996 925
rect 1161 919 1163 931
rect 1200 919 1202 931
rect 1221 919 1223 931
rect 1254 919 1256 931
rect 1275 919 1277 931
rect 1310 919 1312 931
rect 1331 919 1333 931
rect 1364 919 1366 931
rect 1385 919 1387 931
rect 1577 932 1583 933
rect 1577 929 1578 932
rect 1542 927 1546 929
rect 1564 928 1578 929
rect 1582 929 1583 932
rect 1582 928 1591 929
rect 1564 927 1591 928
rect 1597 927 1601 929
rect 1569 922 1575 923
rect 1542 920 1546 922
rect 1564 920 1570 922
rect 993 913 999 914
rect 1569 918 1570 920
rect 1574 919 1575 922
rect 1574 918 1578 919
rect 1569 917 1578 918
rect 1582 917 1591 919
rect 1597 917 1601 919
rect 993 909 994 913
rect 998 909 999 913
rect 993 908 999 909
rect 993 905 995 908
rect 1161 907 1163 913
rect 1200 907 1202 913
rect 1221 907 1223 913
rect 1254 907 1256 913
rect 1275 907 1277 913
rect 1310 907 1312 913
rect 1331 907 1333 913
rect 1364 907 1366 913
rect 1385 907 1387 913
rect 1576 912 1582 913
rect 1576 909 1577 912
rect 1551 907 1555 909
rect 1567 908 1577 909
rect 1581 909 1582 912
rect 1581 908 1591 909
rect 1567 907 1591 908
rect 1597 907 1601 909
rect 974 898 976 902
rect 1612 918 1614 939
rect 1644 936 1646 942
rect 1634 934 1640 935
rect 1644 934 1649 936
rect 1676 934 1680 936
rect 1634 930 1635 934
rect 1639 930 1640 934
rect 1634 928 1640 930
rect 1618 926 1622 928
rect 1631 926 1646 928
rect 1644 920 1646 926
rect 2471 928 2473 932
rect 2478 928 2480 932
rect 2685 930 2687 934
rect 1644 918 1649 920
rect 1667 918 1671 920
rect 1692 919 1696 921
rect 1723 920 1732 921
rect 1723 919 1727 920
rect 1612 916 1622 918
rect 1631 916 1636 918
rect 1640 913 1646 914
rect 1640 910 1641 913
rect 1634 909 1641 910
rect 1645 910 1646 913
rect 1726 916 1727 919
rect 1731 918 1741 920
rect 1753 918 1758 920
rect 2458 919 2460 923
rect 1731 916 1732 918
rect 1726 915 1732 916
rect 1736 911 1741 913
rect 1753 911 1758 913
rect 1645 909 1649 910
rect 1634 908 1649 909
rect 1667 908 1671 910
rect 1701 909 1705 911
rect 1723 910 1738 911
rect 1723 909 1727 910
rect 1614 906 1619 908
rect 1631 906 1636 908
rect 1640 903 1646 904
rect 1640 901 1641 903
rect 1614 899 1619 901
rect 1631 899 1641 901
rect 1645 900 1646 903
rect 1726 906 1727 909
rect 1731 909 1738 910
rect 1731 906 1732 909
rect 1726 905 1732 906
rect 1736 901 1741 903
rect 1750 901 1760 903
rect 1645 899 1649 900
rect 1640 898 1649 899
rect 1676 898 1680 900
rect 1701 899 1705 901
rect 1723 899 1728 901
rect 940 891 942 896
rect 947 891 949 896
rect 907 889 932 891
rect 986 891 988 896
rect 993 891 995 896
rect 1438 888 1440 892
rect 1726 893 1728 899
rect 1726 891 1741 893
rect 1750 891 1754 893
rect 179 869 181 873
rect 189 869 191 873
rect 199 869 201 873
rect 508 871 510 875
rect 518 871 520 875
rect 528 871 530 875
rect 835 874 837 878
rect 845 874 847 878
rect 855 874 857 878
rect 1085 873 1087 875
rect 179 855 181 863
rect 175 854 181 855
rect 189 854 191 863
rect 199 854 201 863
rect 508 857 510 865
rect 175 850 176 854
rect 180 850 181 854
rect 195 853 201 854
rect 175 849 181 850
rect 179 836 181 849
rect 189 847 191 850
rect 195 849 196 853
rect 200 849 201 853
rect 504 856 510 857
rect 518 856 520 865
rect 528 856 530 865
rect 835 860 837 868
rect 504 852 505 856
rect 509 852 510 856
rect 524 855 530 856
rect 504 851 510 852
rect 195 848 201 849
rect 185 846 191 847
rect 185 842 186 846
rect 190 842 191 846
rect 185 841 191 842
rect 186 836 188 841
rect 199 839 201 848
rect 508 838 510 851
rect 518 849 520 852
rect 524 851 525 855
rect 529 851 530 855
rect 831 859 837 860
rect 845 859 847 868
rect 855 859 857 868
rect 1157 873 1159 879
rect 1196 873 1198 879
rect 1217 873 1219 879
rect 1250 873 1252 879
rect 1271 873 1273 879
rect 1306 873 1308 879
rect 1327 873 1329 879
rect 1360 873 1362 879
rect 1381 873 1383 879
rect 1426 877 1428 882
rect 831 855 832 859
rect 836 855 837 859
rect 851 858 857 859
rect 831 854 837 855
rect 524 850 530 851
rect 514 848 520 849
rect 514 844 515 848
rect 519 844 520 848
rect 514 843 520 844
rect 515 838 517 843
rect 528 841 530 850
rect 835 841 837 854
rect 845 852 847 855
rect 851 854 852 858
rect 856 854 857 858
rect 1085 856 1087 867
rect 851 853 857 854
rect 841 851 847 852
rect 841 847 842 851
rect 846 847 847 851
rect 841 846 847 847
rect 842 841 844 846
rect 855 844 857 853
rect 1157 855 1159 867
rect 1196 855 1198 867
rect 1217 855 1219 867
rect 1250 855 1252 867
rect 1271 855 1273 867
rect 1306 855 1308 867
rect 1327 855 1329 867
rect 1360 855 1362 867
rect 1381 855 1383 867
rect 1732 889 1738 891
rect 1732 885 1733 889
rect 1737 885 1738 889
rect 1692 883 1696 885
rect 1723 883 1728 885
rect 1732 884 1738 885
rect 1726 877 1728 883
rect 1758 880 1760 901
rect 1771 910 1775 912
rect 1781 911 1805 912
rect 1781 910 1791 911
rect 1790 907 1791 910
rect 1795 910 1805 911
rect 1817 910 1821 912
rect 1795 907 1796 910
rect 1790 906 1796 907
rect 1771 900 1775 902
rect 1781 900 1790 902
rect 1794 901 1803 902
rect 1794 900 1798 901
rect 1797 897 1798 900
rect 1802 899 1803 901
rect 1802 897 1808 899
rect 1826 897 1830 899
rect 2458 898 2460 907
rect 2471 905 2473 910
rect 2468 904 2474 905
rect 2468 900 2469 904
rect 2473 900 2474 904
rect 2468 899 2474 900
rect 2458 897 2464 898
rect 1797 896 1803 897
rect 2458 893 2459 897
rect 2463 893 2464 897
rect 2468 896 2470 899
rect 2478 897 2480 910
rect 2708 927 2710 947
rect 2715 927 2717 932
rect 2733 930 2735 934
rect 2743 930 2745 934
rect 2753 930 2755 934
rect 2698 918 2700 923
rect 2478 896 2484 897
rect 2458 892 2464 893
rect 2478 892 2479 896
rect 2483 892 2484 896
rect 1771 890 1775 892
rect 1781 891 1808 892
rect 1781 890 1790 891
rect 1789 887 1790 890
rect 1794 890 1808 891
rect 1826 890 1830 892
rect 1794 887 1795 890
rect 1789 886 1795 887
rect 2458 883 2460 892
rect 2468 883 2470 892
rect 2478 891 2484 892
rect 2685 892 2687 905
rect 2698 902 2700 905
rect 2831 930 2833 934
rect 2838 930 2840 934
rect 2818 921 2820 925
rect 2691 901 2700 902
rect 2691 897 2692 901
rect 2696 900 2700 901
rect 2696 897 2697 900
rect 2708 899 2710 902
rect 2691 896 2697 897
rect 2685 891 2691 892
rect 2478 883 2480 891
rect 2685 887 2686 891
rect 2690 887 2691 891
rect 2685 886 2691 887
rect 2685 883 2687 886
rect 2695 883 2697 896
rect 2705 898 2710 899
rect 2705 894 2706 898
rect 2705 893 2710 894
rect 2715 899 2717 902
rect 2733 899 2735 902
rect 2743 899 2745 902
rect 2753 899 2755 902
rect 2818 900 2820 909
rect 2831 907 2833 912
rect 2828 906 2834 907
rect 2828 902 2829 906
rect 2833 902 2834 906
rect 2828 901 2834 902
rect 2818 899 2824 900
rect 2715 898 2737 899
rect 2715 894 2725 898
rect 2729 894 2732 898
rect 2736 894 2737 898
rect 2715 893 2737 894
rect 2741 898 2747 899
rect 2741 894 2742 898
rect 2746 894 2747 898
rect 2741 893 2747 894
rect 2751 898 2757 899
rect 2751 894 2752 898
rect 2756 894 2757 898
rect 2751 893 2757 894
rect 2818 895 2819 899
rect 2823 895 2824 899
rect 2828 898 2830 901
rect 2838 899 2840 912
rect 2838 898 2844 899
rect 2818 894 2824 895
rect 2838 894 2839 898
rect 2843 894 2844 898
rect 2705 890 2707 893
rect 2715 890 2717 893
rect 2735 890 2737 893
rect 2742 890 2744 893
rect 1748 878 1760 880
rect 1748 877 1750 878
rect 1726 875 1736 877
rect 1745 875 1750 877
rect 1726 874 1728 875
rect 1711 873 1728 874
rect 1711 869 1712 873
rect 1716 872 1728 873
rect 1716 869 1717 872
rect 1711 868 1717 869
rect 2458 873 2460 877
rect 2468 873 2470 877
rect 2478 873 2480 877
rect 1655 866 1661 867
rect 1655 863 1656 866
rect 1644 862 1656 863
rect 1660 862 1661 866
rect 2685 866 2687 870
rect 2695 868 2697 873
rect 2705 871 2707 876
rect 2715 871 2717 876
rect 2753 884 2755 893
rect 2818 885 2820 894
rect 2828 885 2830 894
rect 2838 893 2844 894
rect 2838 885 2840 893
rect 2818 875 2820 879
rect 2828 875 2830 879
rect 2838 875 2840 879
rect 2735 866 2737 870
rect 2742 866 2744 870
rect 2753 866 2755 870
rect 1644 861 1661 862
rect 1644 860 1646 861
rect 1426 857 1428 860
rect 1438 857 1440 860
rect 1622 858 1627 860
rect 1636 858 1646 860
rect 1622 857 1624 858
rect 199 823 201 827
rect 528 825 530 829
rect 855 828 857 832
rect 1085 834 1087 852
rect 1197 851 1198 855
rect 1218 851 1219 855
rect 1251 851 1252 855
rect 1272 851 1273 855
rect 1307 851 1308 855
rect 1328 851 1329 855
rect 1361 851 1362 855
rect 1382 851 1383 855
rect 1422 856 1428 857
rect 1422 852 1423 856
rect 1427 852 1428 856
rect 1422 851 1428 852
rect 1434 856 1440 857
rect 1434 852 1435 856
rect 1439 852 1440 856
rect 1434 851 1440 852
rect 1085 828 1087 831
rect 1157 833 1159 851
rect 1196 836 1198 851
rect 1217 836 1219 851
rect 1250 836 1252 851
rect 1271 836 1273 851
rect 1306 836 1308 851
rect 1327 836 1329 851
rect 1360 836 1362 851
rect 1381 836 1383 851
rect 1426 848 1428 851
rect 1438 848 1440 851
rect 1612 855 1624 857
rect 1426 833 1428 838
rect 1612 834 1614 855
rect 1644 852 1646 858
rect 2320 855 2322 860
rect 2327 855 2329 860
rect 2383 860 2408 862
rect 2366 855 2368 860
rect 2373 855 2375 860
rect 1634 850 1640 851
rect 1644 850 1649 852
rect 1676 850 1680 852
rect 1634 846 1635 850
rect 1639 846 1640 850
rect 1634 844 1640 846
rect 2339 849 2341 853
rect 1618 842 1622 844
rect 1631 842 1646 844
rect 1644 836 1646 842
rect 2320 843 2322 846
rect 2316 842 2322 843
rect 2316 838 2317 842
rect 2321 838 2322 842
rect 2316 837 2322 838
rect 1644 834 1649 836
rect 1667 834 1671 836
rect 1157 827 1159 830
rect 1196 827 1198 830
rect 1217 827 1219 830
rect 1250 827 1252 830
rect 1271 827 1273 830
rect 1306 827 1308 830
rect 1327 827 1329 830
rect 1360 827 1362 830
rect 1381 827 1383 830
rect 1438 829 1440 834
rect 1612 832 1622 834
rect 1631 832 1636 834
rect 1640 829 1646 830
rect 1640 826 1641 829
rect 179 814 181 818
rect 186 814 188 818
rect 508 816 510 820
rect 515 816 517 820
rect 835 819 837 823
rect 842 819 844 823
rect 1634 825 1641 826
rect 1645 826 1646 829
rect 2319 826 2321 837
rect 2327 832 2329 846
rect 2383 852 2385 860
rect 2393 852 2395 856
rect 2406 852 2408 860
rect 2467 860 2492 862
rect 2450 855 2452 860
rect 2457 855 2459 860
rect 2406 850 2411 852
rect 2409 847 2411 850
rect 2339 835 2341 843
rect 2335 834 2341 835
rect 2366 834 2368 843
rect 2373 840 2375 843
rect 2373 838 2377 840
rect 2383 838 2385 843
rect 2393 840 2395 843
rect 2393 839 2402 840
rect 2375 834 2377 838
rect 2393 835 2397 839
rect 2401 835 2402 839
rect 2467 852 2469 860
rect 2477 852 2479 856
rect 2490 852 2492 860
rect 2552 855 2554 860
rect 2559 855 2561 860
rect 2680 857 2682 862
rect 2687 857 2689 862
rect 2743 862 2768 864
rect 2726 857 2728 862
rect 2733 857 2735 862
rect 2490 850 2495 852
rect 2493 847 2495 850
rect 2393 834 2402 835
rect 2327 829 2331 832
rect 2335 830 2336 834
rect 2340 830 2341 834
rect 2335 829 2341 830
rect 2329 826 2331 829
rect 2339 826 2341 829
rect 2365 833 2371 834
rect 2365 829 2366 833
rect 2370 829 2371 833
rect 2365 828 2371 829
rect 2375 833 2381 834
rect 2375 829 2376 833
rect 2380 829 2381 833
rect 2393 830 2395 834
rect 2409 830 2411 838
rect 2450 834 2452 843
rect 2457 840 2459 843
rect 2457 838 2461 840
rect 2467 838 2469 843
rect 2477 840 2479 843
rect 2477 839 2486 840
rect 2459 834 2461 838
rect 2477 835 2481 839
rect 2485 835 2486 839
rect 2571 849 2573 853
rect 2552 843 2554 846
rect 2548 842 2554 843
rect 2548 838 2549 842
rect 2553 838 2554 842
rect 2477 834 2486 835
rect 2449 833 2455 834
rect 2375 828 2381 829
rect 2385 828 2395 830
rect 2401 828 2414 830
rect 1645 825 1649 826
rect 1634 824 1649 825
rect 1667 824 1671 826
rect 1614 822 1619 824
rect 1631 822 1636 824
rect 1161 811 1163 814
rect 1200 811 1202 814
rect 1221 811 1223 814
rect 1254 811 1256 814
rect 1275 811 1277 814
rect 1310 811 1312 814
rect 1331 811 1333 814
rect 1364 811 1366 814
rect 1385 811 1387 814
rect 171 802 173 806
rect 95 794 101 795
rect 85 786 87 791
rect 95 790 96 794
rect 100 790 101 794
rect 95 789 101 790
rect 95 784 97 789
rect 105 784 107 789
rect 156 786 162 787
rect 156 782 157 786
rect 161 782 162 786
rect 156 781 162 782
rect 85 771 87 774
rect 95 771 97 774
rect 85 770 91 771
rect 85 766 86 770
rect 90 766 91 770
rect 95 768 99 771
rect 85 765 91 766
rect 85 757 87 765
rect 97 754 99 768
rect 105 763 107 774
rect 160 772 162 781
rect 207 802 209 806
rect 255 802 257 806
rect 187 793 189 797
rect 197 793 199 797
rect 240 786 246 787
rect 240 782 241 786
rect 245 782 246 786
rect 240 781 246 782
rect 171 772 173 775
rect 187 772 189 775
rect 197 772 199 775
rect 207 772 209 775
rect 160 770 173 772
rect 179 770 189 772
rect 193 771 199 772
rect 104 762 110 763
rect 163 762 165 770
rect 179 766 181 770
rect 193 767 194 771
rect 198 767 199 771
rect 193 766 199 767
rect 203 771 209 772
rect 203 767 204 771
rect 208 767 209 771
rect 244 772 246 781
rect 291 802 293 806
rect 271 793 273 797
rect 281 793 283 797
rect 500 804 502 808
rect 424 796 430 797
rect 327 794 333 795
rect 317 786 319 791
rect 327 790 328 794
rect 332 790 333 794
rect 327 789 333 790
rect 255 772 257 775
rect 271 772 273 775
rect 281 772 283 775
rect 291 772 293 775
rect 327 784 329 789
rect 337 784 339 789
rect 414 788 416 793
rect 424 792 425 796
rect 429 792 430 796
rect 424 791 430 792
rect 424 786 426 791
rect 434 786 436 791
rect 485 788 491 789
rect 485 784 486 788
rect 490 784 491 788
rect 485 783 491 784
rect 244 770 257 772
rect 263 770 273 772
rect 277 771 283 772
rect 203 766 209 767
rect 172 765 181 766
rect 104 758 105 762
rect 109 758 110 762
rect 104 757 110 758
rect 104 754 106 757
rect 85 747 87 751
rect 172 761 173 765
rect 177 761 181 765
rect 197 762 199 766
rect 172 760 181 761
rect 179 757 181 760
rect 189 757 191 762
rect 197 760 201 762
rect 199 757 201 760
rect 206 757 208 766
rect 247 762 249 770
rect 263 766 265 770
rect 277 767 278 771
rect 282 767 283 771
rect 277 766 283 767
rect 287 771 293 772
rect 287 767 288 771
rect 292 767 293 771
rect 287 766 293 767
rect 317 771 319 774
rect 327 771 329 774
rect 317 770 323 771
rect 317 766 318 770
rect 322 766 323 770
rect 327 768 331 771
rect 256 765 265 766
rect 163 750 165 753
rect 163 748 168 750
rect 97 740 99 745
rect 104 740 106 745
rect 166 740 168 748
rect 179 744 181 748
rect 189 740 191 748
rect 256 761 257 765
rect 261 761 265 765
rect 281 762 283 766
rect 256 760 265 761
rect 263 757 265 760
rect 273 757 275 762
rect 281 760 285 762
rect 283 757 285 760
rect 290 757 292 766
rect 317 765 323 766
rect 317 757 319 765
rect 247 750 249 753
rect 247 748 252 750
rect 199 740 201 745
rect 206 740 208 745
rect 166 738 191 740
rect 250 740 252 748
rect 263 744 265 748
rect 273 740 275 748
rect 329 754 331 768
rect 337 763 339 774
rect 414 773 416 776
rect 424 773 426 776
rect 414 772 420 773
rect 414 768 415 772
rect 419 768 420 772
rect 424 770 428 773
rect 414 767 420 768
rect 336 762 342 763
rect 336 758 337 762
rect 341 758 342 762
rect 414 759 416 767
rect 336 757 342 758
rect 336 754 338 757
rect 317 747 319 751
rect 426 756 428 770
rect 434 765 436 776
rect 489 774 491 783
rect 536 804 538 808
rect 584 804 586 808
rect 516 795 518 799
rect 526 795 528 799
rect 569 788 575 789
rect 569 784 570 788
rect 574 784 575 788
rect 569 783 575 784
rect 500 774 502 777
rect 516 774 518 777
rect 526 774 528 777
rect 536 774 538 777
rect 489 772 502 774
rect 508 772 518 774
rect 522 773 528 774
rect 433 764 439 765
rect 492 764 494 772
rect 508 768 510 772
rect 522 769 523 773
rect 527 769 528 773
rect 522 768 528 769
rect 532 773 538 774
rect 532 769 533 773
rect 537 769 538 773
rect 573 774 575 783
rect 620 804 622 808
rect 600 795 602 799
rect 610 795 612 799
rect 827 807 829 811
rect 751 799 757 800
rect 656 796 662 797
rect 646 788 648 793
rect 656 792 657 796
rect 661 792 662 796
rect 656 791 662 792
rect 741 791 743 796
rect 751 795 752 799
rect 756 795 757 799
rect 751 794 757 795
rect 584 774 586 777
rect 600 774 602 777
rect 610 774 612 777
rect 620 774 622 777
rect 656 786 658 791
rect 666 786 668 791
rect 751 789 753 794
rect 761 789 763 794
rect 812 791 818 792
rect 812 787 813 791
rect 817 787 818 791
rect 812 786 818 787
rect 741 776 743 779
rect 751 776 753 779
rect 573 772 586 774
rect 592 772 602 774
rect 606 773 612 774
rect 532 768 538 769
rect 501 767 510 768
rect 433 760 434 764
rect 438 760 439 764
rect 433 759 439 760
rect 433 756 435 759
rect 414 749 416 753
rect 501 763 502 767
rect 506 763 510 767
rect 526 764 528 768
rect 501 762 510 763
rect 508 759 510 762
rect 518 759 520 764
rect 526 762 530 764
rect 528 759 530 762
rect 535 759 537 768
rect 576 764 578 772
rect 592 768 594 772
rect 606 769 607 773
rect 611 769 612 773
rect 606 768 612 769
rect 616 773 622 774
rect 616 769 617 773
rect 621 769 622 773
rect 616 768 622 769
rect 646 773 648 776
rect 656 773 658 776
rect 646 772 652 773
rect 646 768 647 772
rect 651 768 652 772
rect 656 770 660 773
rect 585 767 594 768
rect 492 752 494 755
rect 492 750 497 752
rect 283 740 285 745
rect 290 740 292 745
rect 250 738 275 740
rect 329 740 331 745
rect 336 740 338 745
rect 426 742 428 747
rect 433 742 435 747
rect 495 742 497 750
rect 508 746 510 750
rect 518 742 520 750
rect 585 763 586 767
rect 590 763 594 767
rect 610 764 612 768
rect 585 762 594 763
rect 592 759 594 762
rect 602 759 604 764
rect 610 762 614 764
rect 612 759 614 762
rect 619 759 621 768
rect 646 767 652 768
rect 646 759 648 767
rect 576 752 578 755
rect 576 750 581 752
rect 528 742 530 747
rect 535 742 537 747
rect 495 740 520 742
rect 579 742 581 750
rect 592 746 594 750
rect 602 742 604 750
rect 658 756 660 770
rect 666 765 668 776
rect 741 775 747 776
rect 741 771 742 775
rect 746 771 747 775
rect 751 773 755 776
rect 741 770 747 771
rect 665 764 671 765
rect 665 760 666 764
rect 670 760 671 764
rect 741 762 743 770
rect 665 759 671 760
rect 665 756 667 759
rect 753 759 755 773
rect 761 768 763 779
rect 816 777 818 786
rect 863 807 865 811
rect 911 807 913 811
rect 843 798 845 802
rect 853 798 855 802
rect 896 791 902 792
rect 896 787 897 791
rect 901 787 902 791
rect 896 786 902 787
rect 827 777 829 780
rect 843 777 845 780
rect 853 777 855 780
rect 863 777 865 780
rect 816 775 829 777
rect 835 775 845 777
rect 849 776 855 777
rect 760 767 766 768
rect 819 767 821 775
rect 835 771 837 775
rect 849 772 850 776
rect 854 772 855 776
rect 849 771 855 772
rect 859 776 865 777
rect 859 772 860 776
rect 864 772 865 776
rect 900 777 902 786
rect 947 807 949 811
rect 927 798 929 802
rect 937 798 939 802
rect 983 799 989 800
rect 973 791 975 796
rect 983 795 984 799
rect 988 795 989 799
rect 983 794 989 795
rect 911 777 913 780
rect 927 777 929 780
rect 937 777 939 780
rect 947 777 949 780
rect 983 789 985 794
rect 993 789 995 794
rect 1161 790 1163 808
rect 1427 809 1429 814
rect 1439 813 1441 818
rect 1640 819 1646 820
rect 1640 817 1641 819
rect 1614 815 1619 817
rect 1631 815 1641 817
rect 1645 816 1646 819
rect 1645 815 1649 816
rect 1640 814 1649 815
rect 1676 814 1680 816
rect 1200 790 1202 805
rect 1221 790 1223 805
rect 1254 790 1256 805
rect 1275 790 1277 805
rect 1310 790 1312 805
rect 1331 790 1333 805
rect 1364 790 1366 805
rect 1385 790 1387 805
rect 1735 821 1741 822
rect 1735 819 1736 821
rect 1709 817 1714 819
rect 1724 817 1736 819
rect 1740 818 1741 821
rect 1740 817 1744 818
rect 1735 816 1744 817
rect 1753 816 1758 818
rect 1703 812 1709 813
rect 1703 808 1704 812
rect 1708 809 1709 812
rect 2319 811 2321 816
rect 2329 811 2331 816
rect 2365 825 2367 828
rect 2375 825 2377 828
rect 2385 825 2387 828
rect 2401 825 2403 828
rect 1727 809 1744 811
rect 1753 809 1758 811
rect 2325 810 2331 811
rect 1708 808 1714 809
rect 1703 807 1714 808
rect 1724 807 1730 809
rect 1427 796 1429 799
rect 1439 796 1441 799
rect 1423 795 1429 796
rect 1423 791 1424 795
rect 1428 791 1429 795
rect 1423 790 1429 791
rect 1435 795 1441 796
rect 1435 791 1436 795
rect 1440 791 1441 795
rect 1435 790 1441 791
rect 1727 802 1733 803
rect 1727 799 1728 802
rect 1707 797 1712 799
rect 1724 798 1728 799
rect 1732 799 1733 802
rect 2325 806 2326 810
rect 2330 806 2331 810
rect 2339 809 2341 814
rect 2325 805 2331 806
rect 1732 798 1741 799
rect 1724 797 1741 798
rect 1747 797 1751 799
rect 1201 786 1202 790
rect 1222 786 1223 790
rect 1255 786 1256 790
rect 1276 786 1277 790
rect 1311 786 1312 790
rect 1332 786 1333 790
rect 1365 786 1366 790
rect 1386 786 1387 790
rect 1427 787 1429 790
rect 1439 787 1441 790
rect 1621 788 1625 790
rect 1631 789 1648 790
rect 1631 788 1640 789
rect 900 775 913 777
rect 919 775 929 777
rect 933 776 939 777
rect 859 771 865 772
rect 828 770 837 771
rect 760 763 761 767
rect 765 763 766 767
rect 760 762 766 763
rect 760 759 762 762
rect 646 749 648 753
rect 741 752 743 756
rect 828 766 829 770
rect 833 766 837 770
rect 853 767 855 771
rect 828 765 837 766
rect 835 762 837 765
rect 845 762 847 767
rect 853 765 857 767
rect 855 762 857 765
rect 862 762 864 771
rect 903 767 905 775
rect 919 771 921 775
rect 933 772 934 776
rect 938 772 939 776
rect 933 771 939 772
rect 943 776 949 777
rect 943 772 944 776
rect 948 772 949 776
rect 943 771 949 772
rect 973 776 975 779
rect 983 776 985 779
rect 973 775 979 776
rect 973 771 974 775
rect 978 771 979 775
rect 983 773 987 776
rect 912 770 921 771
rect 819 755 821 758
rect 819 753 824 755
rect 612 742 614 747
rect 619 742 621 747
rect 579 740 604 742
rect 658 742 660 747
rect 665 742 667 747
rect 753 745 755 750
rect 760 745 762 750
rect 822 745 824 753
rect 835 749 837 753
rect 845 745 847 753
rect 912 766 913 770
rect 917 766 921 770
rect 937 767 939 771
rect 912 765 921 766
rect 919 762 921 765
rect 929 762 931 767
rect 937 765 941 767
rect 939 762 941 765
rect 946 762 948 771
rect 973 770 979 771
rect 973 762 975 770
rect 903 755 905 758
rect 903 753 908 755
rect 855 745 857 750
rect 862 745 864 750
rect 822 743 847 745
rect 906 745 908 753
rect 919 749 921 753
rect 929 745 931 753
rect 985 759 987 773
rect 993 768 995 779
rect 1161 774 1163 786
rect 1200 774 1202 786
rect 1221 774 1223 786
rect 1254 774 1256 786
rect 1275 774 1277 786
rect 1310 774 1312 786
rect 1331 774 1333 786
rect 1364 774 1366 786
rect 1385 774 1387 786
rect 992 767 998 768
rect 992 763 993 767
rect 997 763 998 767
rect 992 762 998 763
rect 1161 762 1163 768
rect 1200 762 1202 768
rect 1221 762 1223 768
rect 1254 762 1256 768
rect 1275 762 1277 768
rect 1310 762 1312 768
rect 1331 762 1333 768
rect 1364 762 1366 768
rect 1385 762 1387 768
rect 1427 765 1429 770
rect 992 759 994 762
rect 973 752 975 756
rect 1639 785 1640 788
rect 1644 788 1648 789
rect 1660 788 1665 790
rect 1644 785 1645 788
rect 1639 784 1645 785
rect 2375 803 2377 807
rect 2385 803 2387 807
rect 2365 794 2367 798
rect 2412 819 2414 828
rect 2449 829 2450 833
rect 2454 829 2455 833
rect 2449 828 2455 829
rect 2459 833 2465 834
rect 2459 829 2460 833
rect 2464 829 2465 833
rect 2477 830 2479 834
rect 2493 830 2495 838
rect 2548 837 2554 838
rect 2459 828 2465 829
rect 2469 828 2479 830
rect 2485 828 2498 830
rect 2449 825 2451 828
rect 2459 825 2461 828
rect 2469 825 2471 828
rect 2485 825 2487 828
rect 2412 818 2418 819
rect 2412 814 2413 818
rect 2417 814 2418 818
rect 2412 813 2418 814
rect 2459 803 2461 807
rect 2469 803 2471 807
rect 2401 794 2403 798
rect 2449 794 2451 798
rect 2496 819 2498 828
rect 2551 826 2553 837
rect 2559 832 2561 846
rect 2699 851 2701 855
rect 2680 845 2682 848
rect 2676 844 2682 845
rect 2571 835 2573 843
rect 2676 840 2677 844
rect 2681 840 2682 844
rect 2676 839 2682 840
rect 2567 834 2573 835
rect 2559 829 2563 832
rect 2567 830 2568 834
rect 2572 830 2573 834
rect 2567 829 2573 830
rect 2561 826 2563 829
rect 2571 826 2573 829
rect 2679 828 2681 839
rect 2687 834 2689 848
rect 2743 854 2745 862
rect 2753 854 2755 858
rect 2766 854 2768 862
rect 2827 862 2852 864
rect 2810 857 2812 862
rect 2817 857 2819 862
rect 2766 852 2771 854
rect 2769 849 2771 852
rect 2699 837 2701 845
rect 2695 836 2701 837
rect 2726 836 2728 845
rect 2733 842 2735 845
rect 2733 840 2737 842
rect 2743 840 2745 845
rect 2753 842 2755 845
rect 2753 841 2762 842
rect 2735 836 2737 840
rect 2753 837 2757 841
rect 2761 837 2762 841
rect 2827 854 2829 862
rect 2837 854 2839 858
rect 2850 854 2852 862
rect 2912 857 2914 862
rect 2919 857 2921 862
rect 2850 852 2855 854
rect 2853 849 2855 852
rect 2753 836 2762 837
rect 2687 831 2691 834
rect 2695 832 2696 836
rect 2700 832 2701 836
rect 2695 831 2701 832
rect 2689 828 2691 831
rect 2699 828 2701 831
rect 2725 835 2731 836
rect 2725 831 2726 835
rect 2730 831 2731 835
rect 2725 830 2731 831
rect 2735 835 2741 836
rect 2735 831 2736 835
rect 2740 831 2741 835
rect 2753 832 2755 836
rect 2769 832 2771 840
rect 2810 836 2812 845
rect 2817 842 2819 845
rect 2817 840 2821 842
rect 2827 840 2829 845
rect 2837 842 2839 845
rect 2837 841 2846 842
rect 2819 836 2821 840
rect 2837 837 2841 841
rect 2845 837 2846 841
rect 2931 851 2933 855
rect 2912 845 2914 848
rect 2908 844 2914 845
rect 2908 840 2909 844
rect 2913 840 2914 844
rect 2837 836 2846 837
rect 2809 835 2815 836
rect 2735 830 2741 831
rect 2745 830 2755 832
rect 2761 830 2774 832
rect 2496 818 2502 819
rect 2496 814 2497 818
rect 2501 814 2502 818
rect 2496 813 2502 814
rect 2551 811 2553 816
rect 2561 811 2563 816
rect 2557 810 2563 811
rect 2557 806 2558 810
rect 2562 806 2563 810
rect 2571 809 2573 814
rect 2679 813 2681 818
rect 2689 813 2691 818
rect 2725 827 2727 830
rect 2735 827 2737 830
rect 2745 827 2747 830
rect 2761 827 2763 830
rect 2685 812 2691 813
rect 2685 808 2686 812
rect 2690 808 2691 812
rect 2699 811 2701 816
rect 2685 807 2691 808
rect 2557 805 2563 806
rect 2485 794 2487 798
rect 2735 805 2737 809
rect 2745 805 2747 809
rect 2725 796 2727 800
rect 2772 821 2774 830
rect 2809 831 2810 835
rect 2814 831 2815 835
rect 2809 830 2815 831
rect 2819 835 2825 836
rect 2819 831 2820 835
rect 2824 831 2825 835
rect 2837 832 2839 836
rect 2853 832 2855 840
rect 2908 839 2914 840
rect 2819 830 2825 831
rect 2829 830 2839 832
rect 2845 830 2858 832
rect 2809 827 2811 830
rect 2819 827 2821 830
rect 2829 827 2831 830
rect 2845 827 2847 830
rect 2772 820 2778 821
rect 2772 816 2773 820
rect 2777 816 2778 820
rect 2772 815 2778 816
rect 2819 805 2821 809
rect 2829 805 2831 809
rect 2761 796 2763 800
rect 2809 796 2811 800
rect 2856 821 2858 830
rect 2911 828 2913 839
rect 2919 834 2921 848
rect 2931 837 2933 845
rect 2927 836 2933 837
rect 2919 831 2923 834
rect 2927 832 2928 836
rect 2932 832 2933 836
rect 2927 831 2933 832
rect 2921 828 2923 831
rect 2931 828 2933 831
rect 2856 820 2862 821
rect 2856 816 2857 820
rect 2861 816 2862 820
rect 2856 815 2862 816
rect 2911 813 2913 818
rect 2921 813 2923 818
rect 2917 812 2923 813
rect 2917 808 2918 812
rect 2922 808 2923 812
rect 2931 811 2933 816
rect 2917 807 2923 808
rect 2845 796 2847 800
rect 2078 786 2080 790
rect 1642 778 1648 780
rect 1658 779 1669 780
rect 1658 778 1664 779
rect 1614 776 1619 778
rect 1628 776 1645 778
rect 1663 775 1664 778
rect 1668 775 1669 779
rect 1663 774 1669 775
rect 1614 769 1619 771
rect 1628 770 1637 771
rect 1628 769 1632 770
rect 1631 766 1632 769
rect 1636 768 1648 770
rect 1658 768 1663 770
rect 1636 766 1637 768
rect 1631 765 1637 766
rect 2002 778 2008 779
rect 1992 770 1994 775
rect 2002 774 2003 778
rect 2007 774 2008 778
rect 2002 773 2008 774
rect 1439 755 1441 759
rect 2002 768 2004 773
rect 2012 768 2014 773
rect 2063 770 2069 771
rect 2063 766 2064 770
rect 2068 766 2069 770
rect 2063 765 2069 766
rect 1992 755 1994 758
rect 2002 755 2004 758
rect 1992 754 1998 755
rect 939 745 941 750
rect 946 745 948 750
rect 906 743 931 745
rect 985 745 987 750
rect 992 745 994 750
rect 1438 748 1440 752
rect 1992 750 1993 754
rect 1997 750 1998 754
rect 2002 752 2006 755
rect 1992 749 1998 750
rect 1426 737 1428 742
rect 178 723 180 727
rect 188 723 190 727
rect 198 723 200 727
rect 507 725 509 729
rect 517 725 519 729
rect 527 725 529 729
rect 834 728 836 732
rect 844 728 846 732
rect 854 728 856 732
rect 1084 731 1086 733
rect 1156 731 1158 737
rect 1195 731 1197 737
rect 1216 731 1218 737
rect 1249 731 1251 737
rect 1270 731 1272 737
rect 1305 731 1307 737
rect 1326 731 1328 737
rect 1359 731 1361 737
rect 1380 731 1382 737
rect 178 709 180 717
rect 174 708 180 709
rect 188 708 190 717
rect 198 708 200 717
rect 507 711 509 719
rect 174 704 175 708
rect 179 704 180 708
rect 194 707 200 708
rect 174 703 180 704
rect 178 690 180 703
rect 188 701 190 704
rect 194 703 195 707
rect 199 703 200 707
rect 503 710 509 711
rect 517 710 519 719
rect 527 710 529 719
rect 834 714 836 722
rect 503 706 504 710
rect 508 706 509 710
rect 523 709 529 710
rect 503 705 509 706
rect 194 702 200 703
rect 184 700 190 701
rect 184 696 185 700
rect 189 696 190 700
rect 184 695 190 696
rect 185 690 187 695
rect 198 693 200 702
rect 507 692 509 705
rect 517 703 519 706
rect 523 705 524 709
rect 528 705 529 709
rect 830 713 836 714
rect 844 713 846 722
rect 854 713 856 722
rect 1084 714 1086 725
rect 830 709 831 713
rect 835 709 836 713
rect 850 712 856 713
rect 830 708 836 709
rect 523 704 529 705
rect 513 702 519 703
rect 513 698 514 702
rect 518 698 519 702
rect 513 697 519 698
rect 514 692 516 697
rect 527 695 529 704
rect 834 695 836 708
rect 844 706 846 709
rect 850 708 851 712
rect 855 708 856 712
rect 1156 713 1158 725
rect 1195 713 1197 725
rect 1216 713 1218 725
rect 1249 713 1251 725
rect 1270 713 1272 725
rect 1305 713 1307 725
rect 1326 713 1328 725
rect 1359 713 1361 725
rect 1380 713 1382 725
rect 1992 741 1994 749
rect 2004 738 2006 752
rect 2012 747 2014 758
rect 2067 756 2069 765
rect 2114 786 2116 790
rect 2162 786 2164 790
rect 2094 777 2096 781
rect 2104 777 2106 781
rect 2147 770 2153 771
rect 2147 766 2148 770
rect 2152 766 2153 770
rect 2147 765 2153 766
rect 2078 756 2080 759
rect 2094 756 2096 759
rect 2104 756 2106 759
rect 2114 756 2116 759
rect 2067 754 2080 756
rect 2086 754 2096 756
rect 2100 755 2106 756
rect 2011 746 2017 747
rect 2070 746 2072 754
rect 2086 750 2088 754
rect 2100 751 2101 755
rect 2105 751 2106 755
rect 2100 750 2106 751
rect 2110 755 2116 756
rect 2110 751 2111 755
rect 2115 751 2116 755
rect 2151 756 2153 765
rect 2198 786 2200 790
rect 2178 777 2180 781
rect 2188 777 2190 781
rect 2234 778 2240 779
rect 2224 770 2226 775
rect 2234 774 2235 778
rect 2239 774 2240 778
rect 2434 778 2436 782
rect 2234 773 2240 774
rect 2162 756 2164 759
rect 2178 756 2180 759
rect 2188 756 2190 759
rect 2198 756 2200 759
rect 2234 768 2236 773
rect 2244 768 2246 773
rect 2358 770 2364 771
rect 2348 762 2350 767
rect 2358 766 2359 770
rect 2363 766 2364 770
rect 2358 765 2364 766
rect 2151 754 2164 756
rect 2170 754 2180 756
rect 2184 755 2190 756
rect 2110 750 2116 751
rect 2079 749 2088 750
rect 2011 742 2012 746
rect 2016 742 2017 746
rect 2011 741 2017 742
rect 2011 738 2013 741
rect 1992 731 1994 735
rect 2079 745 2080 749
rect 2084 745 2088 749
rect 2104 746 2106 750
rect 2079 744 2088 745
rect 2086 741 2088 744
rect 2096 741 2098 746
rect 2104 744 2108 746
rect 2106 741 2108 744
rect 2113 741 2115 750
rect 2154 746 2156 754
rect 2170 750 2172 754
rect 2184 751 2185 755
rect 2189 751 2190 755
rect 2184 750 2190 751
rect 2194 755 2200 756
rect 2194 751 2195 755
rect 2199 751 2200 755
rect 2194 750 2200 751
rect 2224 755 2226 758
rect 2234 755 2236 758
rect 2224 754 2230 755
rect 2224 750 2225 754
rect 2229 750 2230 754
rect 2234 752 2238 755
rect 2163 749 2172 750
rect 2070 734 2072 737
rect 2070 732 2075 734
rect 2004 724 2006 729
rect 2011 724 2013 729
rect 2073 724 2075 732
rect 2086 728 2088 732
rect 2096 724 2098 732
rect 2163 745 2164 749
rect 2168 745 2172 749
rect 2188 746 2190 750
rect 2163 744 2172 745
rect 2170 741 2172 744
rect 2180 741 2182 746
rect 2188 744 2192 746
rect 2190 741 2192 744
rect 2197 741 2199 750
rect 2224 749 2230 750
rect 2224 741 2226 749
rect 2154 734 2156 737
rect 2154 732 2159 734
rect 2106 724 2108 729
rect 2113 724 2115 729
rect 2073 722 2098 724
rect 2157 724 2159 732
rect 2170 728 2172 732
rect 2180 724 2182 732
rect 2236 738 2238 752
rect 2244 747 2246 758
rect 2358 760 2360 765
rect 2368 760 2370 765
rect 2419 762 2425 763
rect 2419 758 2420 762
rect 2424 758 2425 762
rect 2419 757 2425 758
rect 2348 747 2350 750
rect 2358 747 2360 750
rect 2243 746 2249 747
rect 2243 742 2244 746
rect 2248 742 2249 746
rect 2243 741 2249 742
rect 2348 746 2354 747
rect 2348 742 2349 746
rect 2353 742 2354 746
rect 2358 744 2362 747
rect 2348 741 2354 742
rect 2243 738 2245 741
rect 2224 731 2226 735
rect 2348 733 2350 741
rect 2190 724 2192 729
rect 2197 724 2199 729
rect 2157 722 2182 724
rect 2236 724 2238 729
rect 2243 724 2245 729
rect 2360 730 2362 744
rect 2368 739 2370 750
rect 2423 748 2425 757
rect 2470 778 2472 782
rect 2518 778 2520 782
rect 2450 769 2452 773
rect 2460 769 2462 773
rect 2503 762 2509 763
rect 2503 758 2504 762
rect 2508 758 2509 762
rect 2503 757 2509 758
rect 2434 748 2436 751
rect 2450 748 2452 751
rect 2460 748 2462 751
rect 2470 748 2472 751
rect 2423 746 2436 748
rect 2442 746 2452 748
rect 2456 747 2462 748
rect 2367 738 2373 739
rect 2426 738 2428 746
rect 2442 742 2444 746
rect 2456 743 2457 747
rect 2461 743 2462 747
rect 2456 742 2462 743
rect 2466 747 2472 748
rect 2466 743 2467 747
rect 2471 743 2472 747
rect 2507 748 2509 757
rect 2554 778 2556 782
rect 2534 769 2536 773
rect 2544 769 2546 773
rect 2794 780 2796 784
rect 2718 772 2724 773
rect 2590 770 2596 771
rect 2580 762 2582 767
rect 2590 766 2591 770
rect 2595 766 2596 770
rect 2590 765 2596 766
rect 2518 748 2520 751
rect 2534 748 2536 751
rect 2544 748 2546 751
rect 2554 748 2556 751
rect 2590 760 2592 765
rect 2600 760 2602 765
rect 2708 764 2710 769
rect 2718 768 2719 772
rect 2723 768 2724 772
rect 2718 767 2724 768
rect 2718 762 2720 767
rect 2728 762 2730 767
rect 2779 764 2785 765
rect 2779 760 2780 764
rect 2784 760 2785 764
rect 2779 759 2785 760
rect 2507 746 2520 748
rect 2526 746 2536 748
rect 2540 747 2546 748
rect 2466 742 2472 743
rect 2435 741 2444 742
rect 2367 734 2368 738
rect 2372 734 2373 738
rect 2367 733 2373 734
rect 2367 730 2369 733
rect 2348 723 2350 727
rect 2435 737 2436 741
rect 2440 737 2444 741
rect 2460 738 2462 742
rect 2435 736 2444 737
rect 2442 733 2444 736
rect 2452 733 2454 738
rect 2460 736 2464 738
rect 2462 733 2464 736
rect 2469 733 2471 742
rect 2510 738 2512 746
rect 2526 742 2528 746
rect 2540 743 2541 747
rect 2545 743 2546 747
rect 2540 742 2546 743
rect 2550 747 2556 748
rect 2550 743 2551 747
rect 2555 743 2556 747
rect 2550 742 2556 743
rect 2580 747 2582 750
rect 2590 747 2592 750
rect 2580 746 2586 747
rect 2580 742 2581 746
rect 2585 742 2586 746
rect 2590 744 2594 747
rect 2519 741 2528 742
rect 2426 726 2428 729
rect 2426 724 2431 726
rect 1426 717 1428 720
rect 1438 717 1440 720
rect 1989 717 1991 721
rect 2000 717 2002 721
rect 2007 717 2009 721
rect 850 707 856 708
rect 840 705 846 706
rect 840 701 841 705
rect 845 701 846 705
rect 840 700 846 701
rect 841 695 843 700
rect 854 698 856 707
rect 198 677 200 681
rect 527 679 529 683
rect 1084 692 1086 710
rect 1196 709 1197 713
rect 1217 709 1218 713
rect 1250 709 1251 713
rect 1271 709 1272 713
rect 1306 709 1307 713
rect 1327 709 1328 713
rect 1360 709 1361 713
rect 1381 709 1382 713
rect 1422 716 1428 717
rect 1422 712 1423 716
rect 1427 712 1428 716
rect 1422 711 1428 712
rect 1434 716 1440 717
rect 1434 712 1435 716
rect 1439 712 1440 716
rect 1434 711 1440 712
rect 1084 686 1086 689
rect 1156 691 1158 709
rect 1195 694 1197 709
rect 1216 694 1218 709
rect 1249 694 1251 709
rect 1270 694 1272 709
rect 1305 694 1307 709
rect 1326 694 1328 709
rect 1359 694 1361 709
rect 1380 694 1382 709
rect 1426 708 1428 711
rect 1438 708 1440 711
rect 1426 693 1428 698
rect 854 682 856 686
rect 1156 685 1158 688
rect 1195 685 1197 688
rect 1216 685 1218 688
rect 1249 685 1251 688
rect 1270 685 1272 688
rect 1305 685 1307 688
rect 1326 685 1328 688
rect 1359 685 1361 688
rect 1380 685 1382 688
rect 1438 689 1440 694
rect 1737 693 1743 694
rect 1737 691 1738 693
rect 1711 689 1716 691
rect 1726 689 1738 691
rect 1742 690 1743 693
rect 1989 694 1991 703
rect 2027 711 2029 716
rect 2037 711 2039 716
rect 2047 714 2049 719
rect 2057 717 2059 721
rect 2360 716 2362 721
rect 2367 716 2369 721
rect 2429 716 2431 724
rect 2442 720 2444 724
rect 2452 716 2454 724
rect 2519 737 2520 741
rect 2524 737 2528 741
rect 2544 738 2546 742
rect 2519 736 2528 737
rect 2526 733 2528 736
rect 2536 733 2538 738
rect 2544 736 2548 738
rect 2546 733 2548 736
rect 2553 733 2555 742
rect 2580 741 2586 742
rect 2580 733 2582 741
rect 2510 726 2512 729
rect 2510 724 2515 726
rect 2462 716 2464 721
rect 2469 716 2471 721
rect 2429 714 2454 716
rect 2513 716 2515 724
rect 2526 720 2528 724
rect 2536 716 2538 724
rect 2592 730 2594 744
rect 2600 739 2602 750
rect 2708 749 2710 752
rect 2718 749 2720 752
rect 2708 748 2714 749
rect 2708 744 2709 748
rect 2713 744 2714 748
rect 2718 746 2722 749
rect 2708 743 2714 744
rect 2599 738 2605 739
rect 2599 734 2600 738
rect 2604 734 2605 738
rect 2708 735 2710 743
rect 2599 733 2605 734
rect 2599 730 2601 733
rect 2580 723 2582 727
rect 2720 732 2722 746
rect 2728 741 2730 752
rect 2783 750 2785 759
rect 2830 780 2832 784
rect 2878 780 2880 784
rect 2810 771 2812 775
rect 2820 771 2822 775
rect 2863 764 2869 765
rect 2863 760 2864 764
rect 2868 760 2869 764
rect 2863 759 2869 760
rect 2794 750 2796 753
rect 2810 750 2812 753
rect 2820 750 2822 753
rect 2830 750 2832 753
rect 2783 748 2796 750
rect 2802 748 2812 750
rect 2816 749 2822 750
rect 2727 740 2733 741
rect 2786 740 2788 748
rect 2802 744 2804 748
rect 2816 745 2817 749
rect 2821 745 2822 749
rect 2816 744 2822 745
rect 2826 749 2832 750
rect 2826 745 2827 749
rect 2831 745 2832 749
rect 2867 750 2869 759
rect 2914 780 2916 784
rect 2894 771 2896 775
rect 2904 771 2906 775
rect 2950 772 2956 773
rect 2940 764 2942 769
rect 2950 768 2951 772
rect 2955 768 2956 772
rect 2950 767 2956 768
rect 2878 750 2880 753
rect 2894 750 2896 753
rect 2904 750 2906 753
rect 2914 750 2916 753
rect 2950 762 2952 767
rect 2960 762 2962 767
rect 2867 748 2880 750
rect 2886 748 2896 750
rect 2900 749 2906 750
rect 2826 744 2832 745
rect 2795 743 2804 744
rect 2727 736 2728 740
rect 2732 736 2733 740
rect 2727 735 2733 736
rect 2727 732 2729 735
rect 2708 725 2710 729
rect 2795 739 2796 743
rect 2800 739 2804 743
rect 2820 740 2822 744
rect 2795 738 2804 739
rect 2802 735 2804 738
rect 2812 735 2814 740
rect 2820 738 2824 740
rect 2822 735 2824 738
rect 2829 735 2831 744
rect 2870 740 2872 748
rect 2886 744 2888 748
rect 2900 745 2901 749
rect 2905 745 2906 749
rect 2900 744 2906 745
rect 2910 749 2916 750
rect 2910 745 2911 749
rect 2915 745 2916 749
rect 2910 744 2916 745
rect 2940 749 2942 752
rect 2950 749 2952 752
rect 2940 748 2946 749
rect 2940 744 2941 748
rect 2945 744 2946 748
rect 2950 746 2954 749
rect 2879 743 2888 744
rect 2786 728 2788 731
rect 2786 726 2791 728
rect 2546 716 2548 721
rect 2553 716 2555 721
rect 2513 714 2538 716
rect 2592 716 2594 721
rect 2599 716 2601 721
rect 2720 718 2722 723
rect 2727 718 2729 723
rect 2789 718 2791 726
rect 2802 722 2804 726
rect 2812 718 2814 726
rect 2879 739 2880 743
rect 2884 739 2888 743
rect 2904 740 2906 744
rect 2879 738 2888 739
rect 2886 735 2888 738
rect 2896 735 2898 740
rect 2904 738 2908 740
rect 2906 735 2908 738
rect 2913 735 2915 744
rect 2940 743 2946 744
rect 2940 735 2942 743
rect 2870 728 2872 731
rect 2870 726 2875 728
rect 2822 718 2824 723
rect 2829 718 2831 723
rect 2789 716 2814 718
rect 2873 718 2875 726
rect 2886 722 2888 726
rect 2896 718 2898 726
rect 2952 732 2954 746
rect 2960 741 2962 752
rect 2959 740 2965 741
rect 2959 736 2960 740
rect 2964 736 2965 740
rect 2959 735 2965 736
rect 2959 732 2961 735
rect 2940 725 2942 729
rect 2906 718 2908 723
rect 2913 718 2915 723
rect 2873 716 2898 718
rect 2952 718 2954 723
rect 2959 718 2961 723
rect 2085 707 2087 711
rect 2095 707 2097 711
rect 2105 707 2107 711
rect 2000 694 2002 697
rect 2007 694 2009 697
rect 2027 694 2029 697
rect 2037 694 2039 697
rect 1987 693 1993 694
rect 1742 689 1746 690
rect 1737 688 1746 689
rect 1755 688 1760 690
rect 1987 689 1988 693
rect 1992 689 1993 693
rect 1987 688 1993 689
rect 1997 693 2003 694
rect 1997 689 1998 693
rect 2002 689 2003 693
rect 1997 688 2003 689
rect 2007 693 2029 694
rect 2007 689 2008 693
rect 2012 689 2015 693
rect 2019 689 2029 693
rect 2007 688 2029 689
rect 2033 693 2039 694
rect 2033 689 2034 693
rect 2038 689 2039 693
rect 2033 688 2039 689
rect 2047 691 2049 704
rect 2057 701 2059 704
rect 2053 700 2059 701
rect 2053 696 2054 700
rect 2058 696 2059 700
rect 2053 695 2059 696
rect 2047 690 2053 691
rect 178 668 180 672
rect 185 668 187 672
rect 507 670 509 674
rect 514 670 516 674
rect 834 673 836 677
rect 841 673 843 677
rect 1705 684 1711 685
rect 1705 680 1706 684
rect 1710 681 1711 684
rect 1989 685 1991 688
rect 1999 685 2001 688
rect 2009 685 2011 688
rect 2022 685 2024 688
rect 2027 685 2029 688
rect 2034 685 2036 688
rect 2047 687 2048 690
rect 2044 686 2048 687
rect 2052 686 2053 690
rect 2044 685 2053 686
rect 1729 681 1746 683
rect 1755 681 1760 683
rect 1710 680 1716 681
rect 1705 679 1716 680
rect 1726 679 1732 681
rect 1160 669 1162 672
rect 1199 669 1201 672
rect 1220 669 1222 672
rect 1253 669 1255 672
rect 1274 669 1276 672
rect 1309 669 1311 672
rect 1330 669 1332 672
rect 1363 669 1365 672
rect 1384 669 1386 672
rect 379 645 381 649
rect 389 647 391 652
rect 399 647 401 652
rect 472 645 474 649
rect 482 647 484 652
rect 492 647 494 652
rect 379 623 381 627
rect 389 623 391 634
rect 399 631 401 634
rect 399 630 405 631
rect 399 626 400 630
rect 404 626 405 630
rect 559 645 561 649
rect 569 647 571 652
rect 579 647 581 652
rect 1160 648 1162 666
rect 1199 648 1201 663
rect 1220 648 1222 663
rect 1253 648 1255 663
rect 1274 648 1276 663
rect 1309 648 1311 663
rect 1330 648 1332 663
rect 1363 648 1365 663
rect 1384 648 1386 663
rect 1729 674 1735 675
rect 1729 671 1730 674
rect 1709 669 1714 671
rect 1726 670 1730 671
rect 1734 671 1735 674
rect 1734 670 1743 671
rect 1726 669 1743 670
rect 1749 669 1753 671
rect 1623 660 1627 662
rect 1633 661 1650 662
rect 1633 660 1642 661
rect 1641 657 1642 660
rect 1646 660 1650 661
rect 1662 660 1667 662
rect 1646 657 1647 660
rect 1641 656 1647 657
rect 2044 682 2046 685
rect 2057 682 2059 695
rect 2085 693 2087 701
rect 2081 692 2087 693
rect 2095 692 2097 701
rect 2105 692 2107 701
rect 2441 699 2443 703
rect 2451 699 2453 703
rect 2461 699 2463 703
rect 2801 701 2803 705
rect 2811 701 2813 705
rect 2821 701 2823 705
rect 2081 688 2082 692
rect 2086 688 2087 692
rect 2101 691 2107 692
rect 2081 687 2087 688
rect 2044 664 2046 669
rect 2085 674 2087 687
rect 2095 685 2097 688
rect 2101 687 2102 691
rect 2106 687 2107 691
rect 2101 686 2107 687
rect 2091 684 2097 685
rect 2091 680 2092 684
rect 2096 680 2097 684
rect 2091 679 2097 680
rect 2092 674 2094 679
rect 2105 677 2107 686
rect 2441 685 2443 693
rect 2437 684 2443 685
rect 2451 684 2453 693
rect 2461 684 2463 693
rect 2801 687 2803 695
rect 2437 680 2438 684
rect 2442 680 2443 684
rect 2457 683 2463 684
rect 2437 679 2443 680
rect 1989 655 1991 657
rect 1999 655 2001 657
rect 1644 650 1650 652
rect 1660 651 1671 652
rect 1660 650 1666 651
rect 1616 648 1621 650
rect 1630 648 1647 650
rect 399 625 405 626
rect 379 622 385 623
rect 379 618 380 622
rect 384 618 385 622
rect 379 617 385 618
rect 389 622 395 623
rect 389 618 390 622
rect 394 618 395 622
rect 389 617 395 618
rect 379 612 381 617
rect 392 612 394 617
rect 399 612 401 625
rect 472 623 474 627
rect 482 623 484 634
rect 492 631 494 634
rect 492 630 498 631
rect 492 626 493 630
rect 497 626 498 630
rect 1200 644 1201 648
rect 1221 644 1222 648
rect 1254 644 1255 648
rect 1275 644 1276 648
rect 1310 644 1311 648
rect 1331 644 1332 648
rect 1364 644 1365 648
rect 1385 644 1386 648
rect 492 625 498 626
rect 472 622 478 623
rect 472 618 473 622
rect 477 618 478 622
rect 472 617 478 618
rect 482 622 488 623
rect 482 618 483 622
rect 487 618 488 622
rect 482 617 488 618
rect 472 612 474 617
rect 485 612 487 617
rect 492 612 494 625
rect 559 623 561 627
rect 569 623 571 634
rect 579 631 581 634
rect 1160 632 1162 644
rect 1199 632 1201 644
rect 1220 632 1222 644
rect 1253 632 1255 644
rect 1274 632 1276 644
rect 1309 632 1311 644
rect 1330 632 1332 644
rect 1363 632 1365 644
rect 1384 632 1386 644
rect 1665 647 1666 650
rect 1670 647 1671 651
rect 1665 646 1671 647
rect 1616 641 1621 643
rect 1630 642 1639 643
rect 1630 641 1634 642
rect 1633 638 1634 641
rect 1638 640 1650 642
rect 1660 640 1665 642
rect 1638 638 1639 640
rect 1633 637 1639 638
rect 1694 643 1698 645
rect 1725 644 1734 645
rect 1725 643 1729 644
rect 1728 640 1729 643
rect 1733 642 1743 644
rect 1755 642 1760 644
rect 1733 640 1734 642
rect 1728 639 1734 640
rect 2009 639 2011 657
rect 2022 655 2024 657
rect 2027 655 2029 657
rect 1738 635 1743 637
rect 1755 635 1760 637
rect 2034 637 2036 657
rect 2057 653 2059 657
rect 2441 666 2443 679
rect 2451 677 2453 680
rect 2457 679 2458 683
rect 2462 679 2463 683
rect 2797 686 2803 687
rect 2811 686 2813 695
rect 2821 686 2823 695
rect 2797 682 2798 686
rect 2802 682 2803 686
rect 2817 685 2823 686
rect 2797 681 2803 682
rect 2457 678 2463 679
rect 2447 676 2453 677
rect 2447 672 2448 676
rect 2452 672 2453 676
rect 2447 671 2453 672
rect 2448 666 2450 671
rect 2461 669 2463 678
rect 2105 661 2107 665
rect 2085 652 2087 656
rect 2092 652 2094 656
rect 2801 668 2803 681
rect 2811 679 2813 682
rect 2817 681 2818 685
rect 2822 681 2823 685
rect 2817 680 2823 681
rect 2807 678 2813 679
rect 2807 674 2808 678
rect 2812 674 2813 678
rect 2807 673 2813 674
rect 2808 668 2810 673
rect 2821 671 2823 680
rect 2461 653 2463 657
rect 2821 655 2823 659
rect 2441 644 2443 648
rect 2448 644 2450 648
rect 2801 646 2803 650
rect 2808 646 2810 650
rect 1703 633 1707 635
rect 1725 634 1740 635
rect 1725 633 1729 634
rect 579 630 585 631
rect 579 626 580 630
rect 584 626 585 630
rect 1728 630 1729 633
rect 1733 633 1740 634
rect 1733 630 1734 633
rect 1728 629 1734 630
rect 579 625 585 626
rect 559 622 565 623
rect 559 618 560 622
rect 564 618 565 622
rect 559 617 565 618
rect 569 622 575 623
rect 569 618 570 622
rect 574 618 575 622
rect 569 617 575 618
rect 559 612 561 617
rect 572 612 574 617
rect 579 612 581 625
rect 1160 620 1162 626
rect 1199 620 1201 626
rect 1220 620 1222 626
rect 1253 620 1255 626
rect 1274 620 1276 626
rect 1309 620 1311 626
rect 1330 620 1332 626
rect 1363 620 1365 626
rect 1384 620 1386 626
rect 1738 625 1743 627
rect 1752 625 1762 627
rect 1703 623 1707 625
rect 1725 623 1730 625
rect 1728 617 1730 623
rect 1728 615 1743 617
rect 1752 615 1756 617
rect 379 599 381 603
rect 392 596 394 601
rect 399 596 401 601
rect 472 599 474 603
rect 485 596 487 601
rect 492 596 494 601
rect 559 599 561 603
rect 1734 613 1740 615
rect 1734 609 1735 613
rect 1739 609 1740 613
rect 1694 607 1698 609
rect 1725 607 1730 609
rect 1734 608 1740 609
rect 572 596 574 601
rect 579 596 581 601
rect 1728 601 1730 607
rect 1760 604 1762 625
rect 1750 602 1762 604
rect 1750 601 1752 602
rect 1728 599 1738 601
rect 1747 599 1752 601
rect 1728 598 1730 599
rect 1713 597 1730 598
rect 1713 593 1714 597
rect 1718 596 1730 597
rect 1718 593 1719 596
rect 1713 592 1719 593
rect 1657 590 1663 591
rect 1657 587 1658 590
rect 1646 586 1658 587
rect 1662 586 1663 590
rect 1646 585 1663 586
rect 1646 584 1648 585
rect 1624 582 1629 584
rect 1638 582 1648 584
rect 1624 581 1626 582
rect 1614 579 1626 581
rect 1579 572 1585 573
rect 1579 569 1580 572
rect 1544 567 1548 569
rect 1566 568 1580 569
rect 1584 569 1585 572
rect 1584 568 1593 569
rect 1566 567 1593 568
rect 1599 567 1603 569
rect 1571 562 1577 563
rect 1544 560 1548 562
rect 1566 560 1572 562
rect 1571 558 1572 560
rect 1576 559 1577 562
rect 1576 558 1580 559
rect 1571 557 1580 558
rect 1584 557 1593 559
rect 1599 557 1603 559
rect 1578 552 1584 553
rect 1578 549 1579 552
rect 1553 547 1557 549
rect 1569 548 1579 549
rect 1583 549 1584 552
rect 1583 548 1593 549
rect 1569 547 1593 548
rect 1599 547 1603 549
rect 1614 558 1616 579
rect 1646 576 1648 582
rect 1636 574 1642 575
rect 1646 574 1651 576
rect 1678 574 1682 576
rect 1636 570 1637 574
rect 1641 570 1642 574
rect 1636 568 1642 570
rect 1620 566 1624 568
rect 1633 566 1648 568
rect 1646 560 1648 566
rect 1646 558 1651 560
rect 1669 558 1673 560
rect 1694 559 1698 561
rect 1725 560 1734 561
rect 1725 559 1729 560
rect 1614 556 1624 558
rect 1633 556 1638 558
rect 1642 553 1648 554
rect 1642 550 1643 553
rect 1636 549 1643 550
rect 1647 550 1648 553
rect 1728 556 1729 559
rect 1733 558 1743 560
rect 1755 558 1760 560
rect 1733 556 1734 558
rect 1728 555 1734 556
rect 1738 551 1743 553
rect 1755 551 1760 553
rect 1647 549 1651 550
rect 1636 548 1651 549
rect 1669 548 1673 550
rect 1703 549 1707 551
rect 1725 550 1740 551
rect 1725 549 1729 550
rect 1616 546 1621 548
rect 1633 546 1638 548
rect 1642 543 1648 544
rect 1642 541 1643 543
rect 1616 539 1621 541
rect 1633 539 1643 541
rect 1647 540 1648 543
rect 1728 546 1729 549
rect 1733 549 1740 550
rect 1733 546 1734 549
rect 1728 545 1734 546
rect 1738 541 1743 543
rect 1752 541 1762 543
rect 1647 539 1651 540
rect 1642 538 1651 539
rect 1678 538 1682 540
rect 1703 539 1707 541
rect 1725 539 1730 541
rect 1728 533 1730 539
rect 1728 531 1743 533
rect 1752 531 1756 533
rect 175 514 177 519
rect 182 514 184 519
rect 195 512 197 516
rect 262 514 264 519
rect 269 514 271 519
rect 282 512 284 516
rect 355 514 357 519
rect 362 514 364 519
rect 375 512 377 516
rect 595 514 597 518
rect 608 516 610 521
rect 615 516 617 521
rect 688 514 690 518
rect 701 516 703 521
rect 708 516 710 521
rect 1734 529 1740 531
rect 1734 525 1735 529
rect 1739 525 1740 529
rect 1694 523 1698 525
rect 1725 523 1730 525
rect 1734 524 1740 525
rect 775 514 777 518
rect 788 516 790 521
rect 795 516 797 521
rect 1728 517 1730 523
rect 1760 520 1762 541
rect 1773 550 1777 552
rect 1783 551 1807 552
rect 1783 550 1793 551
rect 1792 547 1793 550
rect 1797 550 1807 551
rect 1819 550 1823 552
rect 1797 547 1798 550
rect 1792 546 1798 547
rect 1773 540 1777 542
rect 1783 540 1792 542
rect 1796 541 1805 542
rect 1796 540 1800 541
rect 1799 537 1800 540
rect 1804 539 1805 541
rect 1804 537 1810 539
rect 1828 537 1832 539
rect 1799 536 1805 537
rect 1773 530 1777 532
rect 1783 531 1810 532
rect 1783 530 1792 531
rect 1791 527 1792 530
rect 1796 530 1810 531
rect 1828 530 1832 532
rect 1796 527 1797 530
rect 1791 526 1797 527
rect 1750 518 1762 520
rect 1750 517 1752 518
rect 1728 515 1738 517
rect 1747 515 1752 517
rect 1728 514 1730 515
rect 1713 513 1730 514
rect 1106 507 1108 509
rect 175 490 177 503
rect 182 498 184 503
rect 195 498 197 503
rect 181 497 187 498
rect 181 493 182 497
rect 186 493 187 497
rect 181 492 187 493
rect 191 497 197 498
rect 191 493 192 497
rect 196 493 197 497
rect 191 492 197 493
rect 171 489 177 490
rect 171 485 172 489
rect 176 485 177 489
rect 171 484 177 485
rect 175 481 177 484
rect 185 481 187 492
rect 195 488 197 492
rect 262 490 264 503
rect 269 498 271 503
rect 282 498 284 503
rect 268 497 274 498
rect 268 493 269 497
rect 273 493 274 497
rect 268 492 274 493
rect 278 497 284 498
rect 278 493 279 497
rect 283 493 284 497
rect 278 492 284 493
rect 258 489 264 490
rect 258 485 259 489
rect 263 485 264 489
rect 258 484 264 485
rect 262 481 264 484
rect 272 481 274 492
rect 282 488 284 492
rect 355 490 357 503
rect 362 498 364 503
rect 375 498 377 503
rect 361 497 367 498
rect 361 493 362 497
rect 366 493 367 497
rect 361 492 367 493
rect 371 497 377 498
rect 371 493 372 497
rect 376 493 377 497
rect 371 492 377 493
rect 351 489 357 490
rect 175 463 177 468
rect 185 463 187 468
rect 195 466 197 470
rect 351 485 352 489
rect 356 485 357 489
rect 351 484 357 485
rect 355 481 357 484
rect 365 481 367 492
rect 375 488 377 492
rect 595 500 597 505
rect 608 500 610 505
rect 595 499 601 500
rect 595 495 596 499
rect 600 495 601 499
rect 595 494 601 495
rect 605 499 611 500
rect 605 495 606 499
rect 610 495 611 499
rect 605 494 611 495
rect 595 490 597 494
rect 262 463 264 468
rect 272 463 274 468
rect 282 466 284 470
rect 605 483 607 494
rect 615 492 617 505
rect 688 500 690 505
rect 701 500 703 505
rect 688 499 694 500
rect 688 495 689 499
rect 693 495 694 499
rect 688 494 694 495
rect 698 499 704 500
rect 698 495 699 499
rect 703 495 704 499
rect 698 494 704 495
rect 615 491 621 492
rect 615 487 616 491
rect 620 487 621 491
rect 688 490 690 494
rect 615 486 621 487
rect 615 483 617 486
rect 355 463 357 468
rect 365 463 367 468
rect 375 466 377 470
rect 595 468 597 472
rect 698 483 700 494
rect 708 492 710 505
rect 775 500 777 505
rect 788 500 790 505
rect 775 499 781 500
rect 775 495 776 499
rect 780 495 781 499
rect 775 494 781 495
rect 785 499 791 500
rect 785 495 786 499
rect 790 495 791 499
rect 785 494 791 495
rect 708 491 714 492
rect 708 487 709 491
rect 713 487 714 491
rect 775 490 777 494
rect 708 486 714 487
rect 708 483 710 486
rect 605 465 607 470
rect 615 465 617 470
rect 688 468 690 472
rect 785 483 787 494
rect 795 492 797 505
rect 1178 507 1180 513
rect 1217 507 1219 513
rect 1238 507 1240 513
rect 1271 507 1273 513
rect 1292 507 1294 513
rect 1327 507 1329 513
rect 1348 507 1350 513
rect 1381 507 1383 513
rect 1402 507 1404 513
rect 1713 509 1714 513
rect 1718 512 1730 513
rect 1718 509 1719 512
rect 1713 508 1719 509
rect 795 491 801 492
rect 795 487 796 491
rect 800 487 801 491
rect 1106 490 1108 501
rect 795 486 801 487
rect 1178 489 1180 501
rect 1217 489 1219 501
rect 1238 489 1240 501
rect 1271 489 1273 501
rect 1292 489 1294 501
rect 1327 489 1329 501
rect 1348 489 1350 501
rect 1381 489 1383 501
rect 1402 489 1404 501
rect 1657 506 1663 507
rect 1657 503 1658 506
rect 1646 502 1658 503
rect 1662 502 1663 506
rect 1646 501 1663 502
rect 1646 500 1648 501
rect 1624 498 1629 500
rect 1638 498 1648 500
rect 1624 497 1626 498
rect 795 483 797 486
rect 698 465 700 470
rect 708 465 710 470
rect 775 468 777 472
rect 785 465 787 470
rect 795 465 797 470
rect 1106 468 1108 486
rect 1218 485 1219 489
rect 1239 485 1240 489
rect 1272 485 1273 489
rect 1293 485 1294 489
rect 1328 485 1329 489
rect 1349 485 1350 489
rect 1382 485 1383 489
rect 1403 485 1404 489
rect 1106 462 1108 465
rect 1178 467 1180 485
rect 1217 470 1219 485
rect 1238 470 1240 485
rect 1271 470 1273 485
rect 1292 470 1294 485
rect 1327 470 1329 485
rect 1348 470 1350 485
rect 1381 470 1383 485
rect 1402 470 1404 485
rect 1614 495 1626 497
rect 1614 474 1616 495
rect 1646 492 1648 498
rect 1636 490 1642 491
rect 1646 490 1651 492
rect 1678 490 1682 492
rect 1636 486 1637 490
rect 1641 486 1642 490
rect 1636 484 1642 486
rect 1620 482 1624 484
rect 1633 482 1648 484
rect 1646 476 1648 482
rect 1646 474 1651 476
rect 1669 474 1673 476
rect 1614 472 1624 474
rect 1633 472 1638 474
rect 1642 469 1648 470
rect 1642 466 1643 469
rect 1636 465 1643 466
rect 1647 466 1648 469
rect 1647 465 1651 466
rect 1636 464 1651 465
rect 1669 464 1673 466
rect 1178 461 1180 464
rect 1217 461 1219 464
rect 1238 461 1240 464
rect 1271 461 1273 464
rect 1292 461 1294 464
rect 1327 461 1329 464
rect 1348 461 1350 464
rect 1381 461 1383 464
rect 1402 461 1404 464
rect 1616 462 1621 464
rect 1633 462 1638 464
rect 1642 459 1648 460
rect 1642 457 1643 459
rect 1616 455 1621 457
rect 1633 455 1643 457
rect 1647 456 1648 459
rect 1647 455 1651 456
rect 1642 454 1651 455
rect 1678 454 1682 456
rect 183 442 185 446
rect 107 434 113 435
rect 97 426 99 431
rect 107 430 108 434
rect 112 430 113 434
rect 107 429 113 430
rect 107 424 109 429
rect 117 424 119 429
rect 168 426 174 427
rect 168 422 169 426
rect 173 422 174 426
rect 168 421 174 422
rect 97 411 99 414
rect 107 411 109 414
rect 97 410 103 411
rect 97 406 98 410
rect 102 406 103 410
rect 107 408 111 411
rect 97 405 103 406
rect 97 397 99 405
rect 109 394 111 408
rect 117 403 119 414
rect 172 412 174 421
rect 219 442 221 446
rect 267 442 269 446
rect 199 433 201 437
rect 209 433 211 437
rect 252 426 258 427
rect 252 422 253 426
rect 257 422 258 426
rect 252 421 258 422
rect 183 412 185 415
rect 199 412 201 415
rect 209 412 211 415
rect 219 412 221 415
rect 172 410 185 412
rect 191 410 201 412
rect 205 411 211 412
rect 116 402 122 403
rect 175 402 177 410
rect 191 406 193 410
rect 205 407 206 411
rect 210 407 211 411
rect 205 406 211 407
rect 215 411 221 412
rect 215 407 216 411
rect 220 407 221 411
rect 256 412 258 421
rect 303 442 305 446
rect 283 433 285 437
rect 293 433 295 437
rect 512 444 514 448
rect 436 436 442 437
rect 339 434 345 435
rect 329 426 331 431
rect 339 430 340 434
rect 344 430 345 434
rect 339 429 345 430
rect 267 412 269 415
rect 283 412 285 415
rect 293 412 295 415
rect 303 412 305 415
rect 339 424 341 429
rect 349 424 351 429
rect 426 428 428 433
rect 436 432 437 436
rect 441 432 442 436
rect 436 431 442 432
rect 436 426 438 431
rect 446 426 448 431
rect 497 428 503 429
rect 497 424 498 428
rect 502 424 503 428
rect 497 423 503 424
rect 256 410 269 412
rect 275 410 285 412
rect 289 411 295 412
rect 215 406 221 407
rect 184 405 193 406
rect 116 398 117 402
rect 121 398 122 402
rect 116 397 122 398
rect 116 394 118 397
rect 97 387 99 391
rect 184 401 185 405
rect 189 401 193 405
rect 209 402 211 406
rect 184 400 193 401
rect 191 397 193 400
rect 201 397 203 402
rect 209 400 213 402
rect 211 397 213 400
rect 218 397 220 406
rect 259 402 261 410
rect 275 406 277 410
rect 289 407 290 411
rect 294 407 295 411
rect 289 406 295 407
rect 299 411 305 412
rect 299 407 300 411
rect 304 407 305 411
rect 299 406 305 407
rect 329 411 331 414
rect 339 411 341 414
rect 329 410 335 411
rect 329 406 330 410
rect 334 406 335 410
rect 339 408 343 411
rect 268 405 277 406
rect 175 390 177 393
rect 175 388 180 390
rect 109 380 111 385
rect 116 380 118 385
rect 178 380 180 388
rect 191 384 193 388
rect 201 380 203 388
rect 268 401 269 405
rect 273 401 277 405
rect 293 402 295 406
rect 268 400 277 401
rect 275 397 277 400
rect 285 397 287 402
rect 293 400 297 402
rect 295 397 297 400
rect 302 397 304 406
rect 329 405 335 406
rect 329 397 331 405
rect 259 390 261 393
rect 259 388 264 390
rect 211 380 213 385
rect 218 380 220 385
rect 178 378 203 380
rect 262 380 264 388
rect 275 384 277 388
rect 285 380 287 388
rect 341 394 343 408
rect 349 403 351 414
rect 426 413 428 416
rect 436 413 438 416
rect 426 412 432 413
rect 426 408 427 412
rect 431 408 432 412
rect 436 410 440 413
rect 426 407 432 408
rect 348 402 354 403
rect 348 398 349 402
rect 353 398 354 402
rect 426 399 428 407
rect 348 397 354 398
rect 348 394 350 397
rect 329 387 331 391
rect 438 396 440 410
rect 446 405 448 416
rect 501 414 503 423
rect 548 444 550 448
rect 596 444 598 448
rect 528 435 530 439
rect 538 435 540 439
rect 581 428 587 429
rect 581 424 582 428
rect 586 424 587 428
rect 581 423 587 424
rect 512 414 514 417
rect 528 414 530 417
rect 538 414 540 417
rect 548 414 550 417
rect 501 412 514 414
rect 520 412 530 414
rect 534 413 540 414
rect 445 404 451 405
rect 504 404 506 412
rect 520 408 522 412
rect 534 409 535 413
rect 539 409 540 413
rect 534 408 540 409
rect 544 413 550 414
rect 544 409 545 413
rect 549 409 550 413
rect 585 414 587 423
rect 632 444 634 448
rect 612 435 614 439
rect 622 435 624 439
rect 839 447 841 451
rect 763 439 769 440
rect 668 436 674 437
rect 658 428 660 433
rect 668 432 669 436
rect 673 432 674 436
rect 668 431 674 432
rect 753 431 755 436
rect 763 435 764 439
rect 768 435 769 439
rect 763 434 769 435
rect 596 414 598 417
rect 612 414 614 417
rect 622 414 624 417
rect 632 414 634 417
rect 668 426 670 431
rect 678 426 680 431
rect 763 429 765 434
rect 773 429 775 434
rect 824 431 830 432
rect 824 427 825 431
rect 829 427 830 431
rect 824 426 830 427
rect 753 416 755 419
rect 763 416 765 419
rect 585 412 598 414
rect 604 412 614 414
rect 618 413 624 414
rect 544 408 550 409
rect 513 407 522 408
rect 445 400 446 404
rect 450 400 451 404
rect 445 399 451 400
rect 445 396 447 399
rect 426 389 428 393
rect 513 403 514 407
rect 518 403 522 407
rect 538 404 540 408
rect 513 402 522 403
rect 520 399 522 402
rect 530 399 532 404
rect 538 402 542 404
rect 540 399 542 402
rect 547 399 549 408
rect 588 404 590 412
rect 604 408 606 412
rect 618 409 619 413
rect 623 409 624 413
rect 618 408 624 409
rect 628 413 634 414
rect 628 409 629 413
rect 633 409 634 413
rect 628 408 634 409
rect 658 413 660 416
rect 668 413 670 416
rect 658 412 664 413
rect 658 408 659 412
rect 663 408 664 412
rect 668 410 672 413
rect 597 407 606 408
rect 504 392 506 395
rect 504 390 509 392
rect 295 380 297 385
rect 302 380 304 385
rect 262 378 287 380
rect 341 380 343 385
rect 348 380 350 385
rect 438 382 440 387
rect 445 382 447 387
rect 507 382 509 390
rect 520 386 522 390
rect 530 382 532 390
rect 597 403 598 407
rect 602 403 606 407
rect 622 404 624 408
rect 597 402 606 403
rect 604 399 606 402
rect 614 399 616 404
rect 622 402 626 404
rect 624 399 626 402
rect 631 399 633 408
rect 658 407 664 408
rect 658 399 660 407
rect 588 392 590 395
rect 588 390 593 392
rect 540 382 542 387
rect 547 382 549 387
rect 507 380 532 382
rect 591 382 593 390
rect 604 386 606 390
rect 614 382 616 390
rect 670 396 672 410
rect 678 405 680 416
rect 753 415 759 416
rect 753 411 754 415
rect 758 411 759 415
rect 763 413 767 416
rect 753 410 759 411
rect 677 404 683 405
rect 677 400 678 404
rect 682 400 683 404
rect 753 402 755 410
rect 677 399 683 400
rect 677 396 679 399
rect 765 399 767 413
rect 773 408 775 419
rect 828 417 830 426
rect 875 447 877 451
rect 923 447 925 451
rect 855 438 857 442
rect 865 438 867 442
rect 908 431 914 432
rect 908 427 909 431
rect 913 427 914 431
rect 908 426 914 427
rect 839 417 841 420
rect 855 417 857 420
rect 865 417 867 420
rect 875 417 877 420
rect 828 415 841 417
rect 847 415 857 417
rect 861 416 867 417
rect 772 407 778 408
rect 831 407 833 415
rect 847 411 849 415
rect 861 412 862 416
rect 866 412 867 416
rect 861 411 867 412
rect 871 416 877 417
rect 871 412 872 416
rect 876 412 877 416
rect 912 417 914 426
rect 959 447 961 451
rect 939 438 941 442
rect 949 438 951 442
rect 1182 445 1184 448
rect 1221 445 1223 448
rect 1242 445 1244 448
rect 1275 445 1277 448
rect 1296 445 1298 448
rect 1331 445 1333 448
rect 1352 445 1354 448
rect 1385 445 1387 448
rect 1406 445 1408 448
rect 1737 461 1743 462
rect 1737 459 1738 461
rect 1711 457 1716 459
rect 1726 457 1738 459
rect 1742 458 1743 461
rect 1742 457 1746 458
rect 1737 456 1746 457
rect 1755 456 1760 458
rect 1705 452 1711 453
rect 1705 448 1706 452
rect 1710 449 1711 452
rect 1729 449 1746 451
rect 1755 449 1760 451
rect 1710 448 1716 449
rect 1705 447 1716 448
rect 1726 447 1732 449
rect 995 439 1001 440
rect 985 431 987 436
rect 995 435 996 439
rect 1000 435 1001 439
rect 995 434 1001 435
rect 923 417 925 420
rect 939 417 941 420
rect 949 417 951 420
rect 959 417 961 420
rect 995 429 997 434
rect 1005 429 1007 434
rect 1182 424 1184 442
rect 1221 424 1223 439
rect 1242 424 1244 439
rect 1275 424 1277 439
rect 1296 424 1298 439
rect 1331 424 1333 439
rect 1352 424 1354 439
rect 1385 424 1387 439
rect 1406 424 1408 439
rect 1729 442 1735 443
rect 1729 439 1730 442
rect 1709 437 1714 439
rect 1726 438 1730 439
rect 1734 439 1735 442
rect 2040 443 2042 448
rect 2047 443 2049 448
rect 1734 438 1743 439
rect 1726 437 1743 438
rect 1749 437 1753 439
rect 1623 428 1627 430
rect 1633 429 1650 430
rect 1633 428 1642 429
rect 1222 420 1223 424
rect 1243 420 1244 424
rect 1276 420 1277 424
rect 1297 420 1298 424
rect 1332 420 1333 424
rect 1353 420 1354 424
rect 1386 420 1387 424
rect 1407 420 1408 424
rect 1641 425 1642 428
rect 1646 428 1650 429
rect 1662 428 1667 430
rect 1646 425 1647 428
rect 1641 424 1647 425
rect 2060 441 2062 445
rect 2127 443 2129 448
rect 2134 443 2136 448
rect 2147 441 2149 445
rect 2220 443 2222 448
rect 2227 443 2229 448
rect 2240 441 2242 445
rect 2460 443 2462 447
rect 2473 445 2475 450
rect 2480 445 2482 450
rect 2553 443 2555 447
rect 2566 445 2568 450
rect 2573 445 2575 450
rect 2640 443 2642 447
rect 2653 445 2655 450
rect 2660 445 2662 450
rect 912 415 925 417
rect 931 415 941 417
rect 945 416 951 417
rect 871 411 877 412
rect 840 410 849 411
rect 772 403 773 407
rect 777 403 778 407
rect 772 402 778 403
rect 772 399 774 402
rect 658 389 660 393
rect 753 392 755 396
rect 840 406 841 410
rect 845 406 849 410
rect 865 407 867 411
rect 840 405 849 406
rect 847 402 849 405
rect 857 402 859 407
rect 865 405 869 407
rect 867 402 869 405
rect 874 402 876 411
rect 915 407 917 415
rect 931 411 933 415
rect 945 412 946 416
rect 950 412 951 416
rect 945 411 951 412
rect 955 416 961 417
rect 955 412 956 416
rect 960 412 961 416
rect 955 411 961 412
rect 985 416 987 419
rect 995 416 997 419
rect 985 415 991 416
rect 985 411 986 415
rect 990 411 991 415
rect 995 413 999 416
rect 924 410 933 411
rect 831 395 833 398
rect 831 393 836 395
rect 624 382 626 387
rect 631 382 633 387
rect 591 380 616 382
rect 670 382 672 387
rect 677 382 679 387
rect 765 385 767 390
rect 772 385 774 390
rect 834 385 836 393
rect 847 389 849 393
rect 857 385 859 393
rect 924 406 925 410
rect 929 406 933 410
rect 949 407 951 411
rect 924 405 933 406
rect 931 402 933 405
rect 941 402 943 407
rect 949 405 953 407
rect 951 402 953 405
rect 958 402 960 411
rect 985 410 991 411
rect 985 402 987 410
rect 915 395 917 398
rect 915 393 920 395
rect 867 385 869 390
rect 874 385 876 390
rect 834 383 859 385
rect 918 385 920 393
rect 931 389 933 393
rect 941 385 943 393
rect 997 399 999 413
rect 1005 408 1007 419
rect 1182 408 1184 420
rect 1221 408 1223 420
rect 1242 408 1244 420
rect 1275 408 1277 420
rect 1296 408 1298 420
rect 1331 408 1333 420
rect 1352 408 1354 420
rect 1385 408 1387 420
rect 1406 408 1408 420
rect 1644 418 1650 420
rect 1660 419 1671 420
rect 1660 418 1666 419
rect 1616 416 1621 418
rect 1630 416 1647 418
rect 1665 415 1666 418
rect 1670 415 1671 419
rect 1665 414 1671 415
rect 2040 419 2042 432
rect 2047 427 2049 432
rect 2060 427 2062 432
rect 2046 426 2052 427
rect 2046 422 2047 426
rect 2051 422 2052 426
rect 2046 421 2052 422
rect 2056 426 2062 427
rect 2056 422 2057 426
rect 2061 422 2062 426
rect 2056 421 2062 422
rect 1616 409 1621 411
rect 1630 410 1639 411
rect 1630 409 1634 410
rect 1004 407 1010 408
rect 1004 403 1005 407
rect 1009 403 1010 407
rect 1004 402 1010 403
rect 1633 406 1634 409
rect 1638 408 1650 410
rect 1660 408 1665 410
rect 1638 406 1639 408
rect 1633 405 1639 406
rect 2036 418 2042 419
rect 2036 414 2037 418
rect 2041 414 2042 418
rect 2036 413 2042 414
rect 2040 410 2042 413
rect 2050 410 2052 421
rect 2060 417 2062 421
rect 2127 419 2129 432
rect 2134 427 2136 432
rect 2147 427 2149 432
rect 2133 426 2139 427
rect 2133 422 2134 426
rect 2138 422 2139 426
rect 2133 421 2139 422
rect 2143 426 2149 427
rect 2143 422 2144 426
rect 2148 422 2149 426
rect 2143 421 2149 422
rect 2123 418 2129 419
rect 1004 399 1006 402
rect 985 392 987 396
rect 1182 396 1184 402
rect 1221 396 1223 402
rect 1242 396 1244 402
rect 1275 396 1277 402
rect 1296 396 1298 402
rect 1331 396 1333 402
rect 1352 396 1354 402
rect 1385 396 1387 402
rect 1406 396 1408 402
rect 2123 414 2124 418
rect 2128 414 2129 418
rect 2123 413 2129 414
rect 2127 410 2129 413
rect 2137 410 2139 421
rect 2147 417 2149 421
rect 2220 419 2222 432
rect 2227 427 2229 432
rect 2240 427 2242 432
rect 2226 426 2232 427
rect 2226 422 2227 426
rect 2231 422 2232 426
rect 2226 421 2232 422
rect 2236 426 2242 427
rect 2236 422 2237 426
rect 2241 422 2242 426
rect 2236 421 2242 422
rect 2216 418 2222 419
rect 951 385 953 390
rect 958 385 960 390
rect 918 383 943 385
rect 997 385 999 390
rect 1004 385 1006 390
rect 2040 392 2042 397
rect 2050 392 2052 397
rect 2060 395 2062 399
rect 2216 414 2217 418
rect 2221 414 2222 418
rect 2216 413 2222 414
rect 2220 410 2222 413
rect 2230 410 2232 421
rect 2240 417 2242 421
rect 2460 429 2462 434
rect 2473 429 2475 434
rect 2460 428 2466 429
rect 2460 424 2461 428
rect 2465 424 2466 428
rect 2460 423 2466 424
rect 2470 428 2476 429
rect 2470 424 2471 428
rect 2475 424 2476 428
rect 2470 423 2476 424
rect 2460 419 2462 423
rect 2127 392 2129 397
rect 2137 392 2139 397
rect 2147 395 2149 399
rect 2470 412 2472 423
rect 2480 421 2482 434
rect 2553 429 2555 434
rect 2566 429 2568 434
rect 2553 428 2559 429
rect 2553 424 2554 428
rect 2558 424 2559 428
rect 2553 423 2559 424
rect 2563 428 2569 429
rect 2563 424 2564 428
rect 2568 424 2569 428
rect 2563 423 2569 424
rect 2480 420 2486 421
rect 2480 416 2481 420
rect 2485 416 2486 420
rect 2553 419 2555 423
rect 2480 415 2486 416
rect 2480 412 2482 415
rect 2220 392 2222 397
rect 2230 392 2232 397
rect 2240 395 2242 399
rect 2460 397 2462 401
rect 2563 412 2565 423
rect 2573 421 2575 434
rect 2640 429 2642 434
rect 2653 429 2655 434
rect 2640 428 2646 429
rect 2640 424 2641 428
rect 2645 424 2646 428
rect 2640 423 2646 424
rect 2650 428 2656 429
rect 2650 424 2651 428
rect 2655 424 2656 428
rect 2650 423 2656 424
rect 2573 420 2579 421
rect 2573 416 2574 420
rect 2578 416 2579 420
rect 2640 419 2642 423
rect 2573 415 2579 416
rect 2573 412 2575 415
rect 2470 394 2472 399
rect 2480 394 2482 399
rect 2553 397 2555 401
rect 2650 412 2652 423
rect 2660 421 2662 434
rect 2660 420 2666 421
rect 2660 416 2661 420
rect 2665 416 2666 420
rect 2660 415 2666 416
rect 2660 412 2662 415
rect 2563 394 2565 399
rect 2573 394 2575 399
rect 2640 397 2642 401
rect 2650 394 2652 399
rect 2660 394 2662 399
rect 190 363 192 367
rect 200 363 202 367
rect 210 363 212 367
rect 519 365 521 369
rect 529 365 531 369
rect 539 365 541 369
rect 846 368 848 372
rect 856 368 858 372
rect 866 368 868 372
rect 2048 371 2050 375
rect 1104 362 1106 364
rect 190 349 192 357
rect 186 348 192 349
rect 200 348 202 357
rect 210 348 212 357
rect 519 351 521 359
rect 186 344 187 348
rect 191 344 192 348
rect 206 347 212 348
rect 186 343 192 344
rect 190 330 192 343
rect 200 341 202 344
rect 206 343 207 347
rect 211 343 212 347
rect 515 350 521 351
rect 529 350 531 359
rect 539 350 541 359
rect 846 354 848 362
rect 515 346 516 350
rect 520 346 521 350
rect 535 349 541 350
rect 515 345 521 346
rect 206 342 212 343
rect 196 340 202 341
rect 196 336 197 340
rect 201 336 202 340
rect 196 335 202 336
rect 197 330 199 335
rect 210 333 212 342
rect 519 332 521 345
rect 529 343 531 346
rect 535 345 536 349
rect 540 345 541 349
rect 842 353 848 354
rect 856 353 858 362
rect 866 353 868 362
rect 1176 362 1178 368
rect 1215 362 1217 368
rect 1236 362 1238 368
rect 1269 362 1271 368
rect 1290 362 1292 368
rect 1325 362 1327 368
rect 1346 362 1348 368
rect 1379 362 1381 368
rect 1400 362 1402 368
rect 1972 363 1978 364
rect 842 349 843 353
rect 847 349 848 353
rect 862 352 868 353
rect 842 348 848 349
rect 535 344 541 345
rect 525 342 531 343
rect 525 338 526 342
rect 530 338 531 342
rect 525 337 531 338
rect 526 332 528 337
rect 539 335 541 344
rect 846 335 848 348
rect 856 346 858 349
rect 862 348 863 352
rect 867 348 868 352
rect 862 347 868 348
rect 852 345 858 346
rect 852 341 853 345
rect 857 341 858 345
rect 852 340 858 341
rect 853 335 855 340
rect 866 338 868 347
rect 1104 345 1106 356
rect 1176 344 1178 356
rect 1215 344 1217 356
rect 1236 344 1238 356
rect 1269 344 1271 356
rect 1290 344 1292 356
rect 1325 344 1327 356
rect 1346 344 1348 356
rect 1379 344 1381 356
rect 1400 344 1402 356
rect 1962 355 1964 360
rect 1972 359 1973 363
rect 1977 359 1978 363
rect 1972 358 1978 359
rect 210 317 212 321
rect 539 319 541 323
rect 866 322 868 326
rect 1104 323 1106 341
rect 1216 340 1217 344
rect 1237 340 1238 344
rect 1270 340 1271 344
rect 1291 340 1292 344
rect 1326 340 1327 344
rect 1347 340 1348 344
rect 1380 340 1381 344
rect 1401 340 1402 344
rect 190 308 192 312
rect 197 308 199 312
rect 519 310 521 314
rect 526 310 528 314
rect 846 313 848 317
rect 853 313 855 317
rect 1104 317 1106 320
rect 1176 322 1178 340
rect 1215 325 1217 340
rect 1236 325 1238 340
rect 1269 325 1271 340
rect 1290 325 1292 340
rect 1325 325 1327 340
rect 1346 325 1348 340
rect 1379 325 1381 340
rect 1400 325 1402 340
rect 1458 336 1460 341
rect 1470 340 1472 345
rect 1972 353 1974 358
rect 1982 353 1984 358
rect 2033 355 2039 356
rect 2033 351 2034 355
rect 2038 351 2039 355
rect 2033 350 2039 351
rect 1729 337 1735 338
rect 1729 335 1730 337
rect 1703 333 1708 335
rect 1718 333 1730 335
rect 1734 334 1735 337
rect 1962 340 1964 343
rect 1972 340 1974 343
rect 1962 339 1968 340
rect 1962 335 1963 339
rect 1967 335 1968 339
rect 1972 337 1976 340
rect 1962 334 1968 335
rect 1734 333 1738 334
rect 1729 332 1738 333
rect 1747 332 1752 334
rect 1458 323 1460 326
rect 1470 323 1472 326
rect 1454 322 1460 323
rect 1176 316 1178 319
rect 1215 316 1217 319
rect 1236 316 1238 319
rect 1269 316 1271 319
rect 1290 316 1292 319
rect 1325 316 1327 319
rect 1346 316 1348 319
rect 1379 316 1381 319
rect 1400 316 1402 319
rect 1454 318 1455 322
rect 1459 318 1460 322
rect 1454 317 1460 318
rect 1466 322 1472 323
rect 1466 318 1467 322
rect 1471 318 1472 322
rect 1466 317 1472 318
rect 1458 314 1460 317
rect 1470 314 1472 317
rect 1697 328 1703 329
rect 1697 324 1698 328
rect 1702 325 1703 328
rect 1721 325 1738 327
rect 1747 325 1752 327
rect 1962 326 1964 334
rect 1702 324 1708 325
rect 1697 323 1708 324
rect 1718 323 1724 325
rect 182 296 184 300
rect 106 288 112 289
rect 96 280 98 285
rect 106 284 107 288
rect 111 284 112 288
rect 106 283 112 284
rect 106 278 108 283
rect 116 278 118 283
rect 167 280 173 281
rect 167 276 168 280
rect 172 276 173 280
rect 167 275 173 276
rect 96 265 98 268
rect 106 265 108 268
rect 96 264 102 265
rect 96 260 97 264
rect 101 260 102 264
rect 106 262 110 265
rect 96 259 102 260
rect 96 251 98 259
rect 108 248 110 262
rect 116 257 118 268
rect 171 266 173 275
rect 218 296 220 300
rect 266 296 268 300
rect 198 287 200 291
rect 208 287 210 291
rect 251 280 257 281
rect 251 276 252 280
rect 256 276 257 280
rect 251 275 257 276
rect 182 266 184 269
rect 198 266 200 269
rect 208 266 210 269
rect 218 266 220 269
rect 171 264 184 266
rect 190 264 200 266
rect 204 265 210 266
rect 115 256 121 257
rect 174 256 176 264
rect 190 260 192 264
rect 204 261 205 265
rect 209 261 210 265
rect 204 260 210 261
rect 214 265 220 266
rect 214 261 215 265
rect 219 261 220 265
rect 255 266 257 275
rect 302 296 304 300
rect 282 287 284 291
rect 292 287 294 291
rect 511 298 513 302
rect 435 290 441 291
rect 338 288 344 289
rect 328 280 330 285
rect 338 284 339 288
rect 343 284 344 288
rect 338 283 344 284
rect 266 266 268 269
rect 282 266 284 269
rect 292 266 294 269
rect 302 266 304 269
rect 338 278 340 283
rect 348 278 350 283
rect 425 282 427 287
rect 435 286 436 290
rect 440 286 441 290
rect 435 285 441 286
rect 435 280 437 285
rect 445 280 447 285
rect 496 282 502 283
rect 496 278 497 282
rect 501 278 502 282
rect 496 277 502 278
rect 255 264 268 266
rect 274 264 284 266
rect 288 265 294 266
rect 214 260 220 261
rect 183 259 192 260
rect 115 252 116 256
rect 120 252 121 256
rect 115 251 121 252
rect 115 248 117 251
rect 96 241 98 245
rect 183 255 184 259
rect 188 255 192 259
rect 208 256 210 260
rect 183 254 192 255
rect 190 251 192 254
rect 200 251 202 256
rect 208 254 212 256
rect 210 251 212 254
rect 217 251 219 260
rect 258 256 260 264
rect 274 260 276 264
rect 288 261 289 265
rect 293 261 294 265
rect 288 260 294 261
rect 298 265 304 266
rect 298 261 299 265
rect 303 261 304 265
rect 298 260 304 261
rect 328 265 330 268
rect 338 265 340 268
rect 328 264 334 265
rect 328 260 329 264
rect 333 260 334 264
rect 338 262 342 265
rect 267 259 276 260
rect 174 244 176 247
rect 174 242 179 244
rect 108 234 110 239
rect 115 234 117 239
rect 177 234 179 242
rect 190 238 192 242
rect 200 234 202 242
rect 267 255 268 259
rect 272 255 276 259
rect 292 256 294 260
rect 267 254 276 255
rect 274 251 276 254
rect 284 251 286 256
rect 292 254 296 256
rect 294 251 296 254
rect 301 251 303 260
rect 328 259 334 260
rect 328 251 330 259
rect 258 244 260 247
rect 258 242 263 244
rect 210 234 212 239
rect 217 234 219 239
rect 177 232 202 234
rect 261 234 263 242
rect 274 238 276 242
rect 284 234 286 242
rect 340 248 342 262
rect 348 257 350 268
rect 425 267 427 270
rect 435 267 437 270
rect 425 266 431 267
rect 425 262 426 266
rect 430 262 431 266
rect 435 264 439 267
rect 425 261 431 262
rect 347 256 353 257
rect 347 252 348 256
rect 352 252 353 256
rect 425 253 427 261
rect 347 251 353 252
rect 347 248 349 251
rect 328 241 330 245
rect 437 250 439 264
rect 445 259 447 270
rect 500 268 502 277
rect 547 298 549 302
rect 595 298 597 302
rect 527 289 529 293
rect 537 289 539 293
rect 580 282 586 283
rect 580 278 581 282
rect 585 278 586 282
rect 580 277 586 278
rect 511 268 513 271
rect 527 268 529 271
rect 537 268 539 271
rect 547 268 549 271
rect 500 266 513 268
rect 519 266 529 268
rect 533 267 539 268
rect 444 258 450 259
rect 503 258 505 266
rect 519 262 521 266
rect 533 263 534 267
rect 538 263 539 267
rect 533 262 539 263
rect 543 267 549 268
rect 543 263 544 267
rect 548 263 549 267
rect 584 268 586 277
rect 631 298 633 302
rect 611 289 613 293
rect 621 289 623 293
rect 838 301 840 305
rect 762 293 768 294
rect 667 290 673 291
rect 657 282 659 287
rect 667 286 668 290
rect 672 286 673 290
rect 667 285 673 286
rect 752 285 754 290
rect 762 289 763 293
rect 767 289 768 293
rect 762 288 768 289
rect 595 268 597 271
rect 611 268 613 271
rect 621 268 623 271
rect 631 268 633 271
rect 667 280 669 285
rect 677 280 679 285
rect 762 283 764 288
rect 772 283 774 288
rect 823 285 829 286
rect 823 281 824 285
rect 828 281 829 285
rect 823 280 829 281
rect 752 270 754 273
rect 762 270 764 273
rect 584 266 597 268
rect 603 266 613 268
rect 617 267 623 268
rect 543 262 549 263
rect 512 261 521 262
rect 444 254 445 258
rect 449 254 450 258
rect 444 253 450 254
rect 444 250 446 253
rect 425 243 427 247
rect 512 257 513 261
rect 517 257 521 261
rect 537 258 539 262
rect 512 256 521 257
rect 519 253 521 256
rect 529 253 531 258
rect 537 256 541 258
rect 539 253 541 256
rect 546 253 548 262
rect 587 258 589 266
rect 603 262 605 266
rect 617 263 618 267
rect 622 263 623 267
rect 617 262 623 263
rect 627 267 633 268
rect 627 263 628 267
rect 632 263 633 267
rect 627 262 633 263
rect 657 267 659 270
rect 667 267 669 270
rect 657 266 663 267
rect 657 262 658 266
rect 662 262 663 266
rect 667 264 671 267
rect 596 261 605 262
rect 503 246 505 249
rect 503 244 508 246
rect 294 234 296 239
rect 301 234 303 239
rect 261 232 286 234
rect 340 234 342 239
rect 347 234 349 239
rect 437 236 439 241
rect 444 236 446 241
rect 506 236 508 244
rect 519 240 521 244
rect 529 236 531 244
rect 596 257 597 261
rect 601 257 605 261
rect 621 258 623 262
rect 596 256 605 257
rect 603 253 605 256
rect 613 253 615 258
rect 621 256 625 258
rect 623 253 625 256
rect 630 253 632 262
rect 657 261 663 262
rect 657 253 659 261
rect 587 246 589 249
rect 587 244 592 246
rect 539 236 541 241
rect 546 236 548 241
rect 506 234 531 236
rect 590 236 592 244
rect 603 240 605 244
rect 613 236 615 244
rect 669 250 671 264
rect 677 259 679 270
rect 752 269 758 270
rect 752 265 753 269
rect 757 265 758 269
rect 762 267 766 270
rect 752 264 758 265
rect 676 258 682 259
rect 676 254 677 258
rect 681 254 682 258
rect 752 256 754 264
rect 676 253 682 254
rect 676 250 678 253
rect 764 253 766 267
rect 772 262 774 273
rect 827 271 829 280
rect 874 301 876 305
rect 922 301 924 305
rect 854 292 856 296
rect 864 292 866 296
rect 907 285 913 286
rect 907 281 908 285
rect 912 281 913 285
rect 907 280 913 281
rect 838 271 840 274
rect 854 271 856 274
rect 864 271 866 274
rect 874 271 876 274
rect 827 269 840 271
rect 846 269 856 271
rect 860 270 866 271
rect 771 261 777 262
rect 830 261 832 269
rect 846 265 848 269
rect 860 266 861 270
rect 865 266 866 270
rect 860 265 866 266
rect 870 270 876 271
rect 870 266 871 270
rect 875 266 876 270
rect 911 271 913 280
rect 958 301 960 305
rect 938 292 940 296
rect 948 292 950 296
rect 1180 300 1182 303
rect 1219 300 1221 303
rect 1240 300 1242 303
rect 1273 300 1275 303
rect 1294 300 1296 303
rect 1329 300 1331 303
rect 1350 300 1352 303
rect 1383 300 1385 303
rect 1404 300 1406 303
rect 994 293 1000 294
rect 984 285 986 290
rect 994 289 995 293
rect 999 289 1000 293
rect 994 288 1000 289
rect 922 271 924 274
rect 938 271 940 274
rect 948 271 950 274
rect 958 271 960 274
rect 994 283 996 288
rect 1004 283 1006 288
rect 1180 279 1182 297
rect 1219 279 1221 294
rect 1240 279 1242 294
rect 1273 279 1275 294
rect 1294 279 1296 294
rect 1329 279 1331 294
rect 1350 279 1352 294
rect 1383 279 1385 294
rect 1404 279 1406 294
rect 1458 292 1460 297
rect 1721 318 1727 319
rect 1721 315 1722 318
rect 1701 313 1706 315
rect 1718 314 1722 315
rect 1726 315 1727 318
rect 1974 323 1976 337
rect 1982 332 1984 343
rect 2037 341 2039 350
rect 2084 371 2086 375
rect 2132 371 2134 375
rect 2064 362 2066 366
rect 2074 362 2076 366
rect 2117 355 2123 356
rect 2117 351 2118 355
rect 2122 351 2123 355
rect 2117 350 2123 351
rect 2048 341 2050 344
rect 2064 341 2066 344
rect 2074 341 2076 344
rect 2084 341 2086 344
rect 2037 339 2050 341
rect 2056 339 2066 341
rect 2070 340 2076 341
rect 1981 331 1987 332
rect 2040 331 2042 339
rect 2056 335 2058 339
rect 2070 336 2071 340
rect 2075 336 2076 340
rect 2070 335 2076 336
rect 2080 340 2086 341
rect 2080 336 2081 340
rect 2085 336 2086 340
rect 2121 341 2123 350
rect 2168 371 2170 375
rect 2148 362 2150 366
rect 2158 362 2160 366
rect 2377 373 2379 377
rect 2301 365 2307 366
rect 2204 363 2210 364
rect 2194 355 2196 360
rect 2204 359 2205 363
rect 2209 359 2210 363
rect 2204 358 2210 359
rect 2132 341 2134 344
rect 2148 341 2150 344
rect 2158 341 2160 344
rect 2168 341 2170 344
rect 2204 353 2206 358
rect 2214 353 2216 358
rect 2291 357 2293 362
rect 2301 361 2302 365
rect 2306 361 2307 365
rect 2301 360 2307 361
rect 2301 355 2303 360
rect 2311 355 2313 360
rect 2362 357 2368 358
rect 2362 353 2363 357
rect 2367 353 2368 357
rect 2362 352 2368 353
rect 2121 339 2134 341
rect 2140 339 2150 341
rect 2154 340 2160 341
rect 2080 335 2086 336
rect 2049 334 2058 335
rect 1981 327 1982 331
rect 1986 327 1987 331
rect 1981 326 1987 327
rect 1981 323 1983 326
rect 1962 316 1964 320
rect 1726 314 1735 315
rect 1718 313 1735 314
rect 1741 313 1745 315
rect 2049 330 2050 334
rect 2054 330 2058 334
rect 2074 331 2076 335
rect 2049 329 2058 330
rect 2056 326 2058 329
rect 2066 326 2068 331
rect 2074 329 2078 331
rect 2076 326 2078 329
rect 2083 326 2085 335
rect 2124 331 2126 339
rect 2140 335 2142 339
rect 2154 336 2155 340
rect 2159 336 2160 340
rect 2154 335 2160 336
rect 2164 340 2170 341
rect 2164 336 2165 340
rect 2169 336 2170 340
rect 2164 335 2170 336
rect 2194 340 2196 343
rect 2204 340 2206 343
rect 2194 339 2200 340
rect 2194 335 2195 339
rect 2199 335 2200 339
rect 2204 337 2208 340
rect 2133 334 2142 335
rect 2040 319 2042 322
rect 2040 317 2045 319
rect 1974 309 1976 314
rect 1981 309 1983 314
rect 2043 309 2045 317
rect 2056 313 2058 317
rect 2066 309 2068 317
rect 2133 330 2134 334
rect 2138 330 2142 334
rect 2158 331 2160 335
rect 2133 329 2142 330
rect 2140 326 2142 329
rect 2150 326 2152 331
rect 2158 329 2162 331
rect 2160 326 2162 329
rect 2167 326 2169 335
rect 2194 334 2200 335
rect 2194 326 2196 334
rect 2124 319 2126 322
rect 2124 317 2129 319
rect 2076 309 2078 314
rect 2083 309 2085 314
rect 2043 307 2068 309
rect 2127 309 2129 317
rect 2140 313 2142 317
rect 2150 309 2152 317
rect 2206 323 2208 337
rect 2214 332 2216 343
rect 2291 342 2293 345
rect 2301 342 2303 345
rect 2291 341 2297 342
rect 2291 337 2292 341
rect 2296 337 2297 341
rect 2301 339 2305 342
rect 2291 336 2297 337
rect 2213 331 2219 332
rect 2213 327 2214 331
rect 2218 327 2219 331
rect 2291 328 2293 336
rect 2213 326 2219 327
rect 2213 323 2215 326
rect 2194 316 2196 320
rect 2303 325 2305 339
rect 2311 334 2313 345
rect 2366 343 2368 352
rect 2413 373 2415 377
rect 2461 373 2463 377
rect 2393 364 2395 368
rect 2403 364 2405 368
rect 2446 357 2452 358
rect 2446 353 2447 357
rect 2451 353 2452 357
rect 2446 352 2452 353
rect 2377 343 2379 346
rect 2393 343 2395 346
rect 2403 343 2405 346
rect 2413 343 2415 346
rect 2366 341 2379 343
rect 2385 341 2395 343
rect 2399 342 2405 343
rect 2310 333 2316 334
rect 2369 333 2371 341
rect 2385 337 2387 341
rect 2399 338 2400 342
rect 2404 338 2405 342
rect 2399 337 2405 338
rect 2409 342 2415 343
rect 2409 338 2410 342
rect 2414 338 2415 342
rect 2450 343 2452 352
rect 2497 373 2499 377
rect 2477 364 2479 368
rect 2487 364 2489 368
rect 2704 376 2706 380
rect 2628 368 2634 369
rect 2533 365 2539 366
rect 2523 357 2525 362
rect 2533 361 2534 365
rect 2538 361 2539 365
rect 2533 360 2539 361
rect 2618 360 2620 365
rect 2628 364 2629 368
rect 2633 364 2634 368
rect 2628 363 2634 364
rect 2461 343 2463 346
rect 2477 343 2479 346
rect 2487 343 2489 346
rect 2497 343 2499 346
rect 2533 355 2535 360
rect 2543 355 2545 360
rect 2628 358 2630 363
rect 2638 358 2640 363
rect 2689 360 2695 361
rect 2689 356 2690 360
rect 2694 356 2695 360
rect 2689 355 2695 356
rect 2618 345 2620 348
rect 2628 345 2630 348
rect 2450 341 2463 343
rect 2469 341 2479 343
rect 2483 342 2489 343
rect 2409 337 2415 338
rect 2378 336 2387 337
rect 2310 329 2311 333
rect 2315 329 2316 333
rect 2310 328 2316 329
rect 2310 325 2312 328
rect 2291 318 2293 322
rect 2378 332 2379 336
rect 2383 332 2387 336
rect 2403 333 2405 337
rect 2378 331 2387 332
rect 2385 328 2387 331
rect 2395 328 2397 333
rect 2403 331 2407 333
rect 2405 328 2407 331
rect 2412 328 2414 337
rect 2453 333 2455 341
rect 2469 337 2471 341
rect 2483 338 2484 342
rect 2488 338 2489 342
rect 2483 337 2489 338
rect 2493 342 2499 343
rect 2493 338 2494 342
rect 2498 338 2499 342
rect 2493 337 2499 338
rect 2523 342 2525 345
rect 2533 342 2535 345
rect 2523 341 2529 342
rect 2523 337 2524 341
rect 2528 337 2529 341
rect 2533 339 2537 342
rect 2462 336 2471 337
rect 2369 321 2371 324
rect 2369 319 2374 321
rect 2160 309 2162 314
rect 2167 309 2169 314
rect 2127 307 2152 309
rect 2206 309 2208 314
rect 2213 309 2215 314
rect 2303 311 2305 316
rect 2310 311 2312 316
rect 2372 311 2374 319
rect 2385 315 2387 319
rect 2395 311 2397 319
rect 2462 332 2463 336
rect 2467 332 2471 336
rect 2487 333 2489 337
rect 2462 331 2471 332
rect 2469 328 2471 331
rect 2479 328 2481 333
rect 2487 331 2491 333
rect 2489 328 2491 331
rect 2496 328 2498 337
rect 2523 336 2529 337
rect 2523 328 2525 336
rect 2453 321 2455 324
rect 2453 319 2458 321
rect 2405 311 2407 316
rect 2412 311 2414 316
rect 2372 309 2397 311
rect 2456 311 2458 319
rect 2469 315 2471 319
rect 2479 311 2481 319
rect 2535 325 2537 339
rect 2543 334 2545 345
rect 2618 344 2624 345
rect 2618 340 2619 344
rect 2623 340 2624 344
rect 2628 342 2632 345
rect 2618 339 2624 340
rect 2542 333 2548 334
rect 2542 329 2543 333
rect 2547 329 2548 333
rect 2618 331 2620 339
rect 2542 328 2548 329
rect 2542 325 2544 328
rect 2630 328 2632 342
rect 2638 337 2640 348
rect 2693 346 2695 355
rect 2740 376 2742 380
rect 2788 376 2790 380
rect 2720 367 2722 371
rect 2730 367 2732 371
rect 2773 360 2779 361
rect 2773 356 2774 360
rect 2778 356 2779 360
rect 2773 355 2779 356
rect 2704 346 2706 349
rect 2720 346 2722 349
rect 2730 346 2732 349
rect 2740 346 2742 349
rect 2693 344 2706 346
rect 2712 344 2722 346
rect 2726 345 2732 346
rect 2637 336 2643 337
rect 2696 336 2698 344
rect 2712 340 2714 344
rect 2726 341 2727 345
rect 2731 341 2732 345
rect 2726 340 2732 341
rect 2736 345 2742 346
rect 2736 341 2737 345
rect 2741 341 2742 345
rect 2777 346 2779 355
rect 2824 376 2826 380
rect 2804 367 2806 371
rect 2814 367 2816 371
rect 2860 368 2866 369
rect 2850 360 2852 365
rect 2860 364 2861 368
rect 2865 364 2866 368
rect 2860 363 2866 364
rect 2788 346 2790 349
rect 2804 346 2806 349
rect 2814 346 2816 349
rect 2824 346 2826 349
rect 2860 358 2862 363
rect 2870 358 2872 363
rect 2777 344 2790 346
rect 2796 344 2806 346
rect 2810 345 2816 346
rect 2736 340 2742 341
rect 2705 339 2714 340
rect 2637 332 2638 336
rect 2642 332 2643 336
rect 2637 331 2643 332
rect 2637 328 2639 331
rect 2523 318 2525 322
rect 2618 321 2620 325
rect 2705 335 2706 339
rect 2710 335 2714 339
rect 2730 336 2732 340
rect 2705 334 2714 335
rect 2712 331 2714 334
rect 2722 331 2724 336
rect 2730 334 2734 336
rect 2732 331 2734 334
rect 2739 331 2741 340
rect 2780 336 2782 344
rect 2796 340 2798 344
rect 2810 341 2811 345
rect 2815 341 2816 345
rect 2810 340 2816 341
rect 2820 345 2826 346
rect 2820 341 2821 345
rect 2825 341 2826 345
rect 2820 340 2826 341
rect 2850 345 2852 348
rect 2860 345 2862 348
rect 2850 344 2856 345
rect 2850 340 2851 344
rect 2855 340 2856 344
rect 2860 342 2864 345
rect 2789 339 2798 340
rect 2696 324 2698 327
rect 2696 322 2701 324
rect 2489 311 2491 316
rect 2496 311 2498 316
rect 2456 309 2481 311
rect 2535 311 2537 316
rect 2542 311 2544 316
rect 2630 314 2632 319
rect 2637 314 2639 319
rect 2699 314 2701 322
rect 2712 318 2714 322
rect 2722 314 2724 322
rect 2789 335 2790 339
rect 2794 335 2798 339
rect 2814 336 2816 340
rect 2789 334 2798 335
rect 2796 331 2798 334
rect 2806 331 2808 336
rect 2814 334 2818 336
rect 2816 331 2818 334
rect 2823 331 2825 340
rect 2850 339 2856 340
rect 2850 331 2852 339
rect 2780 324 2782 327
rect 2780 322 2785 324
rect 2732 314 2734 319
rect 2739 314 2741 319
rect 2699 312 2724 314
rect 2783 314 2785 322
rect 2796 318 2798 322
rect 2806 314 2808 322
rect 2862 328 2864 342
rect 2870 337 2872 348
rect 2869 336 2875 337
rect 2869 332 2870 336
rect 2874 332 2875 336
rect 2869 331 2875 332
rect 2869 328 2871 331
rect 2850 321 2852 325
rect 2816 314 2818 319
rect 2823 314 2825 319
rect 2783 312 2808 314
rect 2862 314 2864 319
rect 2869 314 2871 319
rect 2055 292 2057 296
rect 2065 292 2067 296
rect 2075 292 2077 296
rect 2384 294 2386 298
rect 2394 294 2396 298
rect 2404 294 2406 298
rect 2711 297 2713 301
rect 2721 297 2723 301
rect 2731 297 2733 301
rect 1686 287 1690 289
rect 1717 288 1726 289
rect 1717 287 1721 288
rect 1470 282 1472 286
rect 1720 284 1721 287
rect 1725 286 1735 288
rect 1747 286 1752 288
rect 1725 284 1726 286
rect 1720 283 1726 284
rect 1730 279 1735 281
rect 1747 279 1752 281
rect 1220 275 1221 279
rect 1241 275 1242 279
rect 1274 275 1275 279
rect 1295 275 1296 279
rect 1330 275 1331 279
rect 1351 275 1352 279
rect 1384 275 1385 279
rect 1405 275 1406 279
rect 1695 277 1699 279
rect 1717 278 1732 279
rect 1717 277 1721 278
rect 911 269 924 271
rect 930 269 940 271
rect 944 270 950 271
rect 870 265 876 266
rect 839 264 848 265
rect 771 257 772 261
rect 776 257 777 261
rect 771 256 777 257
rect 771 253 773 256
rect 657 243 659 247
rect 752 246 754 250
rect 839 260 840 264
rect 844 260 848 264
rect 864 261 866 265
rect 839 259 848 260
rect 846 256 848 259
rect 856 256 858 261
rect 864 259 868 261
rect 866 256 868 259
rect 873 256 875 265
rect 914 261 916 269
rect 930 265 932 269
rect 944 266 945 270
rect 949 266 950 270
rect 944 265 950 266
rect 954 270 960 271
rect 954 266 955 270
rect 959 266 960 270
rect 954 265 960 266
rect 984 270 986 273
rect 994 270 996 273
rect 984 269 990 270
rect 984 265 985 269
rect 989 265 990 269
rect 994 267 998 270
rect 923 264 932 265
rect 830 249 832 252
rect 830 247 835 249
rect 623 236 625 241
rect 630 236 632 241
rect 590 234 615 236
rect 669 236 671 241
rect 676 236 678 241
rect 764 239 766 244
rect 771 239 773 244
rect 833 239 835 247
rect 846 243 848 247
rect 856 239 858 247
rect 923 260 924 264
rect 928 260 932 264
rect 948 261 950 265
rect 923 259 932 260
rect 930 256 932 259
rect 940 256 942 261
rect 948 259 952 261
rect 950 256 952 259
rect 957 256 959 265
rect 984 264 990 265
rect 984 256 986 264
rect 914 249 916 252
rect 914 247 919 249
rect 866 239 868 244
rect 873 239 875 244
rect 833 237 858 239
rect 917 239 919 247
rect 930 243 932 247
rect 940 239 942 247
rect 996 253 998 267
rect 1004 262 1006 273
rect 1180 263 1182 275
rect 1219 263 1221 275
rect 1240 263 1242 275
rect 1273 263 1275 275
rect 1294 263 1296 275
rect 1329 263 1331 275
rect 1350 263 1352 275
rect 1383 263 1385 275
rect 1404 263 1406 275
rect 1720 274 1721 277
rect 1725 277 1732 278
rect 2055 278 2057 286
rect 1725 274 1726 277
rect 1720 273 1726 274
rect 2051 277 2057 278
rect 2065 277 2067 286
rect 2075 277 2077 286
rect 2384 280 2386 288
rect 2051 273 2052 277
rect 2056 273 2057 277
rect 2071 276 2077 277
rect 2051 272 2057 273
rect 1730 269 1735 271
rect 1744 269 1754 271
rect 1695 267 1699 269
rect 1717 267 1722 269
rect 1003 261 1009 262
rect 1003 257 1004 261
rect 1008 257 1009 261
rect 1720 261 1722 267
rect 1720 259 1735 261
rect 1744 259 1748 261
rect 1003 256 1009 257
rect 1003 253 1005 256
rect 984 246 986 250
rect 1180 251 1182 257
rect 1219 251 1221 257
rect 1240 251 1242 257
rect 1273 251 1275 257
rect 1294 251 1296 257
rect 1329 251 1331 257
rect 1350 251 1352 257
rect 1383 251 1385 257
rect 1404 251 1406 257
rect 1472 253 1474 257
rect 1726 257 1732 259
rect 1726 253 1727 257
rect 1731 253 1732 257
rect 950 239 952 244
rect 957 239 959 244
rect 917 237 942 239
rect 996 239 998 244
rect 1003 239 1005 244
rect 1460 242 1462 247
rect 189 217 191 221
rect 199 217 201 221
rect 209 217 211 221
rect 518 219 520 223
rect 528 219 530 223
rect 538 219 540 223
rect 845 222 847 226
rect 855 222 857 226
rect 865 222 867 226
rect 1105 220 1107 222
rect 189 203 191 211
rect 185 202 191 203
rect 199 202 201 211
rect 209 202 211 211
rect 518 205 520 213
rect 185 198 186 202
rect 190 198 191 202
rect 205 201 211 202
rect 185 197 191 198
rect 189 184 191 197
rect 199 195 201 198
rect 205 197 206 201
rect 210 197 211 201
rect 514 204 520 205
rect 528 204 530 213
rect 538 204 540 213
rect 845 208 847 216
rect 514 200 515 204
rect 519 200 520 204
rect 534 203 540 204
rect 514 199 520 200
rect 205 196 211 197
rect 195 194 201 195
rect 195 190 196 194
rect 200 190 201 194
rect 195 189 201 190
rect 196 184 198 189
rect 209 187 211 196
rect 518 186 520 199
rect 528 197 530 200
rect 534 199 535 203
rect 539 199 540 203
rect 841 207 847 208
rect 855 207 857 216
rect 865 207 867 216
rect 1177 220 1179 226
rect 1216 220 1218 226
rect 1237 220 1239 226
rect 1270 220 1272 226
rect 1291 220 1293 226
rect 1326 220 1328 226
rect 1347 220 1349 226
rect 1380 220 1382 226
rect 1401 220 1403 226
rect 1686 251 1690 253
rect 1717 251 1722 253
rect 1726 252 1732 253
rect 1720 245 1722 251
rect 1752 248 1754 269
rect 2055 259 2057 272
rect 2065 270 2067 273
rect 2071 272 2072 276
rect 2076 272 2077 276
rect 2380 279 2386 280
rect 2394 279 2396 288
rect 2404 279 2406 288
rect 2711 283 2713 291
rect 2380 275 2381 279
rect 2385 275 2386 279
rect 2400 278 2406 279
rect 2380 274 2386 275
rect 2071 271 2077 272
rect 2061 269 2067 270
rect 2061 265 2062 269
rect 2066 265 2067 269
rect 2061 264 2067 265
rect 2062 259 2064 264
rect 2075 262 2077 271
rect 1742 246 1754 248
rect 1742 245 1744 246
rect 1720 243 1730 245
rect 1739 243 1744 245
rect 1720 242 1722 243
rect 1705 241 1722 242
rect 1705 237 1706 241
rect 1710 240 1722 241
rect 1710 237 1711 240
rect 1705 236 1711 237
rect 2384 261 2386 274
rect 2394 272 2396 275
rect 2400 274 2401 278
rect 2405 274 2406 278
rect 2707 282 2713 283
rect 2721 282 2723 291
rect 2731 282 2733 291
rect 2707 278 2708 282
rect 2712 278 2713 282
rect 2727 281 2733 282
rect 2707 277 2713 278
rect 2400 273 2406 274
rect 2390 271 2396 272
rect 2390 267 2391 271
rect 2395 267 2396 271
rect 2390 266 2396 267
rect 2391 261 2393 266
rect 2404 264 2406 273
rect 2711 264 2713 277
rect 2721 275 2723 278
rect 2727 277 2728 281
rect 2732 277 2733 281
rect 2727 276 2733 277
rect 2717 274 2723 275
rect 2717 270 2718 274
rect 2722 270 2723 274
rect 2717 269 2723 270
rect 2718 264 2720 269
rect 2731 267 2733 276
rect 2075 246 2077 250
rect 2404 248 2406 252
rect 2731 251 2733 255
rect 2055 237 2057 241
rect 2062 237 2064 241
rect 2384 239 2386 243
rect 2391 239 2393 243
rect 2711 242 2713 246
rect 2718 242 2720 246
rect 1460 222 1462 225
rect 1472 222 1474 225
rect 2047 225 2049 229
rect 1456 221 1462 222
rect 1456 217 1457 221
rect 1461 217 1462 221
rect 1456 216 1462 217
rect 1468 221 1474 222
rect 1468 217 1469 221
rect 1473 217 1474 221
rect 1468 216 1474 217
rect 841 203 842 207
rect 846 203 847 207
rect 861 206 867 207
rect 841 202 847 203
rect 534 198 540 199
rect 524 196 530 197
rect 524 192 525 196
rect 529 192 530 196
rect 524 191 530 192
rect 525 186 527 191
rect 538 189 540 198
rect 845 189 847 202
rect 855 200 857 203
rect 861 202 862 206
rect 866 202 867 206
rect 1105 203 1107 214
rect 861 201 867 202
rect 851 199 857 200
rect 851 195 852 199
rect 856 195 857 199
rect 851 194 857 195
rect 852 189 854 194
rect 865 192 867 201
rect 1177 202 1179 214
rect 1216 202 1218 214
rect 1237 202 1239 214
rect 1270 202 1272 214
rect 1291 202 1293 214
rect 1326 202 1328 214
rect 1347 202 1349 214
rect 1380 202 1382 214
rect 1401 202 1403 214
rect 1460 213 1462 216
rect 1472 213 1474 216
rect 1971 217 1977 218
rect 209 171 211 175
rect 538 173 540 177
rect 865 176 867 180
rect 1105 181 1107 199
rect 1217 198 1218 202
rect 1238 198 1239 202
rect 1271 198 1272 202
rect 1292 198 1293 202
rect 1327 198 1328 202
rect 1348 198 1349 202
rect 1381 198 1382 202
rect 1402 198 1403 202
rect 1460 198 1462 203
rect 1961 209 1963 214
rect 1971 213 1972 217
rect 1976 213 1977 217
rect 1971 212 1977 213
rect 1686 203 1690 205
rect 1717 204 1726 205
rect 1717 203 1721 204
rect 1105 175 1107 178
rect 1177 180 1179 198
rect 1216 183 1218 198
rect 1237 183 1239 198
rect 1270 183 1272 198
rect 1291 183 1293 198
rect 1326 183 1328 198
rect 1347 183 1349 198
rect 1380 183 1382 198
rect 1401 183 1403 198
rect 1472 194 1474 199
rect 1720 200 1721 203
rect 1725 202 1735 204
rect 1747 202 1752 204
rect 1725 200 1726 202
rect 1720 199 1726 200
rect 1730 195 1735 197
rect 1747 195 1752 197
rect 1695 193 1699 195
rect 1717 194 1732 195
rect 1717 193 1721 194
rect 1720 190 1721 193
rect 1725 193 1732 194
rect 1725 190 1726 193
rect 1720 189 1726 190
rect 1730 185 1735 187
rect 1744 185 1754 187
rect 1695 183 1699 185
rect 1717 183 1722 185
rect 1177 174 1179 177
rect 1216 174 1218 177
rect 1237 174 1239 177
rect 1270 174 1272 177
rect 1291 174 1293 177
rect 1326 174 1328 177
rect 1347 174 1349 177
rect 1380 174 1382 177
rect 1401 174 1403 177
rect 1720 177 1722 183
rect 1720 175 1735 177
rect 1744 175 1748 177
rect 189 162 191 166
rect 196 162 198 166
rect 518 164 520 168
rect 525 164 527 168
rect 845 167 847 171
rect 852 167 854 171
rect 1726 173 1732 175
rect 1726 169 1727 173
rect 1731 169 1732 173
rect 1686 167 1690 169
rect 1717 167 1722 169
rect 1726 168 1732 169
rect 1181 158 1183 161
rect 1220 158 1222 161
rect 1241 158 1243 161
rect 1274 158 1276 161
rect 1295 158 1297 161
rect 1330 158 1332 161
rect 1351 158 1353 161
rect 1384 158 1386 161
rect 1405 158 1407 161
rect 390 139 392 143
rect 400 141 402 146
rect 410 141 412 146
rect 483 139 485 143
rect 493 141 495 146
rect 503 141 505 146
rect 390 117 392 121
rect 400 117 402 128
rect 410 125 412 128
rect 410 124 416 125
rect 410 120 411 124
rect 415 120 416 124
rect 570 139 572 143
rect 580 141 582 146
rect 590 141 592 146
rect 410 119 416 120
rect 390 116 396 117
rect 390 112 391 116
rect 395 112 396 116
rect 390 111 396 112
rect 400 116 406 117
rect 400 112 401 116
rect 405 112 406 116
rect 400 111 406 112
rect 390 106 392 111
rect 403 106 405 111
rect 410 106 412 119
rect 483 117 485 121
rect 493 117 495 128
rect 503 125 505 128
rect 503 124 509 125
rect 503 120 504 124
rect 508 120 509 124
rect 1181 137 1183 155
rect 1462 157 1464 162
rect 1474 161 1476 166
rect 1220 137 1222 152
rect 1241 137 1243 152
rect 1274 137 1276 152
rect 1295 137 1297 152
rect 1330 137 1332 152
rect 1351 137 1353 152
rect 1384 137 1386 152
rect 1405 137 1407 152
rect 1720 161 1722 167
rect 1752 164 1754 185
rect 1971 207 1973 212
rect 1981 207 1983 212
rect 2032 209 2038 210
rect 2032 205 2033 209
rect 2037 205 2038 209
rect 2032 204 2038 205
rect 1765 194 1769 196
rect 1775 195 1799 196
rect 1775 194 1785 195
rect 1784 191 1785 194
rect 1789 194 1799 195
rect 1811 194 1815 196
rect 1961 194 1963 197
rect 1971 194 1973 197
rect 1789 191 1790 194
rect 1784 190 1790 191
rect 1961 193 1967 194
rect 1765 184 1769 186
rect 1775 184 1784 186
rect 1788 185 1797 186
rect 1788 184 1792 185
rect 1791 181 1792 184
rect 1796 183 1797 185
rect 1961 189 1962 193
rect 1966 189 1967 193
rect 1971 191 1975 194
rect 1961 188 1967 189
rect 1796 181 1802 183
rect 1820 181 1824 183
rect 1791 180 1797 181
rect 1961 180 1963 188
rect 1765 174 1769 176
rect 1775 175 1802 176
rect 1775 174 1784 175
rect 1783 171 1784 174
rect 1788 174 1802 175
rect 1820 174 1824 176
rect 1973 177 1975 191
rect 1981 186 1983 197
rect 2036 195 2038 204
rect 2083 225 2085 229
rect 2131 225 2133 229
rect 2063 216 2065 220
rect 2073 216 2075 220
rect 2116 209 2122 210
rect 2116 205 2117 209
rect 2121 205 2122 209
rect 2116 204 2122 205
rect 2047 195 2049 198
rect 2063 195 2065 198
rect 2073 195 2075 198
rect 2083 195 2085 198
rect 2036 193 2049 195
rect 2055 193 2065 195
rect 2069 194 2075 195
rect 1980 185 1986 186
rect 2039 185 2041 193
rect 2055 189 2057 193
rect 2069 190 2070 194
rect 2074 190 2075 194
rect 2069 189 2075 190
rect 2079 194 2085 195
rect 2079 190 2080 194
rect 2084 190 2085 194
rect 2120 195 2122 204
rect 2167 225 2169 229
rect 2147 216 2149 220
rect 2157 216 2159 220
rect 2376 227 2378 231
rect 2300 219 2306 220
rect 2203 217 2209 218
rect 2193 209 2195 214
rect 2203 213 2204 217
rect 2208 213 2209 217
rect 2203 212 2209 213
rect 2131 195 2133 198
rect 2147 195 2149 198
rect 2157 195 2159 198
rect 2167 195 2169 198
rect 2203 207 2205 212
rect 2213 207 2215 212
rect 2290 211 2292 216
rect 2300 215 2301 219
rect 2305 215 2306 219
rect 2300 214 2306 215
rect 2300 209 2302 214
rect 2310 209 2312 214
rect 2361 211 2367 212
rect 2361 207 2362 211
rect 2366 207 2367 211
rect 2361 206 2367 207
rect 2120 193 2133 195
rect 2139 193 2149 195
rect 2153 194 2159 195
rect 2079 189 2085 190
rect 2048 188 2057 189
rect 1980 181 1981 185
rect 1985 181 1986 185
rect 1980 180 1986 181
rect 1980 177 1982 180
rect 1788 171 1789 174
rect 1783 170 1789 171
rect 1961 170 1963 174
rect 2048 184 2049 188
rect 2053 184 2057 188
rect 2073 185 2075 189
rect 2048 183 2057 184
rect 2055 180 2057 183
rect 2065 180 2067 185
rect 2073 183 2077 185
rect 2075 180 2077 183
rect 2082 180 2084 189
rect 2123 185 2125 193
rect 2139 189 2141 193
rect 2153 190 2154 194
rect 2158 190 2159 194
rect 2153 189 2159 190
rect 2163 194 2169 195
rect 2163 190 2164 194
rect 2168 190 2169 194
rect 2163 189 2169 190
rect 2193 194 2195 197
rect 2203 194 2205 197
rect 2193 193 2199 194
rect 2193 189 2194 193
rect 2198 189 2199 193
rect 2203 191 2207 194
rect 2132 188 2141 189
rect 2039 173 2041 176
rect 2039 171 2044 173
rect 1742 162 1754 164
rect 1973 163 1975 168
rect 1980 163 1982 168
rect 2042 163 2044 171
rect 2055 167 2057 171
rect 2065 163 2067 171
rect 2132 184 2133 188
rect 2137 184 2141 188
rect 2157 185 2159 189
rect 2132 183 2141 184
rect 2139 180 2141 183
rect 2149 180 2151 185
rect 2157 183 2161 185
rect 2159 180 2161 183
rect 2166 180 2168 189
rect 2193 188 2199 189
rect 2193 180 2195 188
rect 2123 173 2125 176
rect 2123 171 2128 173
rect 2075 163 2077 168
rect 2082 163 2084 168
rect 1742 161 1744 162
rect 2042 161 2067 163
rect 2126 163 2128 171
rect 2139 167 2141 171
rect 2149 163 2151 171
rect 2205 177 2207 191
rect 2213 186 2215 197
rect 2290 196 2292 199
rect 2300 196 2302 199
rect 2290 195 2296 196
rect 2290 191 2291 195
rect 2295 191 2296 195
rect 2300 193 2304 196
rect 2290 190 2296 191
rect 2212 185 2218 186
rect 2212 181 2213 185
rect 2217 181 2218 185
rect 2290 182 2292 190
rect 2212 180 2218 181
rect 2212 177 2214 180
rect 2193 170 2195 174
rect 2302 179 2304 193
rect 2310 188 2312 199
rect 2365 197 2367 206
rect 2412 227 2414 231
rect 2460 227 2462 231
rect 2392 218 2394 222
rect 2402 218 2404 222
rect 2445 211 2451 212
rect 2445 207 2446 211
rect 2450 207 2451 211
rect 2445 206 2451 207
rect 2376 197 2378 200
rect 2392 197 2394 200
rect 2402 197 2404 200
rect 2412 197 2414 200
rect 2365 195 2378 197
rect 2384 195 2394 197
rect 2398 196 2404 197
rect 2309 187 2315 188
rect 2368 187 2370 195
rect 2384 191 2386 195
rect 2398 192 2399 196
rect 2403 192 2404 196
rect 2398 191 2404 192
rect 2408 196 2414 197
rect 2408 192 2409 196
rect 2413 192 2414 196
rect 2449 197 2451 206
rect 2496 227 2498 231
rect 2476 218 2478 222
rect 2486 218 2488 222
rect 2703 230 2705 234
rect 2627 222 2633 223
rect 2532 219 2538 220
rect 2522 211 2524 216
rect 2532 215 2533 219
rect 2537 215 2538 219
rect 2532 214 2538 215
rect 2617 214 2619 219
rect 2627 218 2628 222
rect 2632 218 2633 222
rect 2627 217 2633 218
rect 2460 197 2462 200
rect 2476 197 2478 200
rect 2486 197 2488 200
rect 2496 197 2498 200
rect 2532 209 2534 214
rect 2542 209 2544 214
rect 2627 212 2629 217
rect 2637 212 2639 217
rect 2688 214 2694 215
rect 2688 210 2689 214
rect 2693 210 2694 214
rect 2688 209 2694 210
rect 2617 199 2619 202
rect 2627 199 2629 202
rect 2449 195 2462 197
rect 2468 195 2478 197
rect 2482 196 2488 197
rect 2408 191 2414 192
rect 2377 190 2386 191
rect 2309 183 2310 187
rect 2314 183 2315 187
rect 2309 182 2315 183
rect 2309 179 2311 182
rect 2290 172 2292 176
rect 2377 186 2378 190
rect 2382 186 2386 190
rect 2402 187 2404 191
rect 2377 185 2386 186
rect 2384 182 2386 185
rect 2394 182 2396 187
rect 2402 185 2406 187
rect 2404 182 2406 185
rect 2411 182 2413 191
rect 2452 187 2454 195
rect 2468 191 2470 195
rect 2482 192 2483 196
rect 2487 192 2488 196
rect 2482 191 2488 192
rect 2492 196 2498 197
rect 2492 192 2493 196
rect 2497 192 2498 196
rect 2492 191 2498 192
rect 2522 196 2524 199
rect 2532 196 2534 199
rect 2522 195 2528 196
rect 2522 191 2523 195
rect 2527 191 2528 195
rect 2532 193 2536 196
rect 2461 190 2470 191
rect 2368 175 2370 178
rect 2368 173 2373 175
rect 2159 163 2161 168
rect 2166 163 2168 168
rect 2126 161 2151 163
rect 2205 163 2207 168
rect 2212 163 2214 168
rect 2302 165 2304 170
rect 2309 165 2311 170
rect 2371 165 2373 173
rect 2384 169 2386 173
rect 2394 165 2396 173
rect 2461 186 2462 190
rect 2466 186 2470 190
rect 2486 187 2488 191
rect 2461 185 2470 186
rect 2468 182 2470 185
rect 2478 182 2480 187
rect 2486 185 2490 187
rect 2488 182 2490 185
rect 2495 182 2497 191
rect 2522 190 2528 191
rect 2522 182 2524 190
rect 2452 175 2454 178
rect 2452 173 2457 175
rect 2404 165 2406 170
rect 2411 165 2413 170
rect 2371 163 2396 165
rect 2455 165 2457 173
rect 2468 169 2470 173
rect 2478 165 2480 173
rect 2534 179 2536 193
rect 2542 188 2544 199
rect 2617 198 2623 199
rect 2617 194 2618 198
rect 2622 194 2623 198
rect 2627 196 2631 199
rect 2617 193 2623 194
rect 2541 187 2547 188
rect 2541 183 2542 187
rect 2546 183 2547 187
rect 2617 185 2619 193
rect 2541 182 2547 183
rect 2541 179 2543 182
rect 2629 182 2631 196
rect 2637 191 2639 202
rect 2692 200 2694 209
rect 2739 230 2741 234
rect 2787 230 2789 234
rect 2719 221 2721 225
rect 2729 221 2731 225
rect 2772 214 2778 215
rect 2772 210 2773 214
rect 2777 210 2778 214
rect 2772 209 2778 210
rect 2703 200 2705 203
rect 2719 200 2721 203
rect 2729 200 2731 203
rect 2739 200 2741 203
rect 2692 198 2705 200
rect 2711 198 2721 200
rect 2725 199 2731 200
rect 2636 190 2642 191
rect 2695 190 2697 198
rect 2711 194 2713 198
rect 2725 195 2726 199
rect 2730 195 2731 199
rect 2725 194 2731 195
rect 2735 199 2741 200
rect 2735 195 2736 199
rect 2740 195 2741 199
rect 2776 200 2778 209
rect 2823 230 2825 234
rect 2803 221 2805 225
rect 2813 221 2815 225
rect 2859 222 2865 223
rect 2849 214 2851 219
rect 2859 218 2860 222
rect 2864 218 2865 222
rect 2859 217 2865 218
rect 2787 200 2789 203
rect 2803 200 2805 203
rect 2813 200 2815 203
rect 2823 200 2825 203
rect 2859 212 2861 217
rect 2869 212 2871 217
rect 2776 198 2789 200
rect 2795 198 2805 200
rect 2809 199 2815 200
rect 2735 194 2741 195
rect 2704 193 2713 194
rect 2636 186 2637 190
rect 2641 186 2642 190
rect 2636 185 2642 186
rect 2636 182 2638 185
rect 2522 172 2524 176
rect 2617 175 2619 179
rect 2704 189 2705 193
rect 2709 189 2713 193
rect 2729 190 2731 194
rect 2704 188 2713 189
rect 2711 185 2713 188
rect 2721 185 2723 190
rect 2729 188 2733 190
rect 2731 185 2733 188
rect 2738 185 2740 194
rect 2779 190 2781 198
rect 2795 194 2797 198
rect 2809 195 2810 199
rect 2814 195 2815 199
rect 2809 194 2815 195
rect 2819 199 2825 200
rect 2819 195 2820 199
rect 2824 195 2825 199
rect 2819 194 2825 195
rect 2849 199 2851 202
rect 2859 199 2861 202
rect 2849 198 2855 199
rect 2849 194 2850 198
rect 2854 194 2855 198
rect 2859 196 2863 199
rect 2788 193 2797 194
rect 2695 178 2697 181
rect 2695 176 2700 178
rect 2488 165 2490 170
rect 2495 165 2497 170
rect 2455 163 2480 165
rect 2534 165 2536 170
rect 2541 165 2543 170
rect 2629 168 2631 173
rect 2636 168 2638 173
rect 2698 168 2700 176
rect 2711 172 2713 176
rect 2721 168 2723 176
rect 2788 189 2789 193
rect 2793 189 2797 193
rect 2813 190 2815 194
rect 2788 188 2797 189
rect 2795 185 2797 188
rect 2805 185 2807 190
rect 2813 188 2817 190
rect 2815 185 2817 188
rect 2822 185 2824 194
rect 2849 193 2855 194
rect 2849 185 2851 193
rect 2779 178 2781 181
rect 2779 176 2784 178
rect 2731 168 2733 173
rect 2738 168 2740 173
rect 2698 166 2723 168
rect 2782 168 2784 176
rect 2795 172 2797 176
rect 2805 168 2807 176
rect 2861 182 2863 196
rect 2869 191 2871 202
rect 2868 190 2874 191
rect 2868 186 2869 190
rect 2873 186 2874 190
rect 2868 185 2874 186
rect 2868 182 2870 185
rect 2849 175 2851 179
rect 2815 168 2817 173
rect 2822 168 2824 173
rect 2782 166 2807 168
rect 2861 168 2863 173
rect 2868 168 2870 173
rect 1720 159 1730 161
rect 1739 159 1744 161
rect 1720 158 1722 159
rect 1705 157 1722 158
rect 1705 153 1706 157
rect 1710 156 1722 157
rect 1710 153 1711 156
rect 1705 152 1711 153
rect 1462 144 1464 147
rect 1474 144 1476 147
rect 1755 146 1759 148
rect 1772 147 1794 148
rect 1772 146 1776 147
rect 1458 143 1464 144
rect 1458 139 1459 143
rect 1463 139 1464 143
rect 1458 138 1464 139
rect 1470 143 1476 144
rect 1470 139 1471 143
rect 1475 139 1476 143
rect 1470 138 1476 139
rect 1775 143 1776 146
rect 1780 146 1794 147
rect 1819 146 1823 148
rect 2054 146 2056 150
rect 2064 146 2066 150
rect 2074 146 2076 150
rect 2383 148 2385 152
rect 2393 148 2395 152
rect 2403 148 2405 152
rect 2710 151 2712 155
rect 2720 151 2722 155
rect 2730 151 2732 155
rect 1780 143 1781 146
rect 1775 142 1781 143
rect 1785 141 1791 142
rect 1785 138 1786 141
rect 1221 133 1222 137
rect 1242 133 1243 137
rect 1275 133 1276 137
rect 1296 133 1297 137
rect 1331 133 1332 137
rect 1352 133 1353 137
rect 1385 133 1386 137
rect 1406 133 1407 137
rect 1462 135 1464 138
rect 1474 135 1476 138
rect 1757 136 1762 138
rect 1772 137 1786 138
rect 1790 137 1791 141
rect 1772 136 1791 137
rect 503 119 509 120
rect 483 116 489 117
rect 483 112 484 116
rect 488 112 489 116
rect 483 111 489 112
rect 493 116 499 117
rect 493 112 494 116
rect 498 112 499 116
rect 493 111 499 112
rect 483 106 485 111
rect 496 106 498 111
rect 503 106 505 119
rect 570 117 572 121
rect 580 117 582 128
rect 590 125 592 128
rect 590 124 596 125
rect 590 120 591 124
rect 595 120 596 124
rect 1181 121 1183 133
rect 1220 121 1222 133
rect 1241 121 1243 133
rect 1274 121 1276 133
rect 1295 121 1297 133
rect 1330 121 1332 133
rect 1351 121 1353 133
rect 1384 121 1386 133
rect 1405 121 1407 133
rect 590 119 596 120
rect 570 116 576 117
rect 570 112 571 116
rect 575 112 576 116
rect 570 111 576 112
rect 580 116 586 117
rect 580 112 581 116
rect 585 112 586 116
rect 580 111 586 112
rect 570 106 572 111
rect 583 106 585 111
rect 590 106 592 119
rect 1181 109 1183 115
rect 1220 109 1222 115
rect 1241 109 1243 115
rect 1274 109 1276 115
rect 1295 109 1297 115
rect 1330 109 1332 115
rect 1351 109 1353 115
rect 1384 109 1386 115
rect 1405 109 1407 115
rect 1462 113 1464 118
rect 390 93 392 97
rect 403 90 405 95
rect 410 90 412 95
rect 483 93 485 97
rect 496 90 498 95
rect 503 90 505 95
rect 570 93 572 97
rect 1789 135 1791 136
rect 1789 133 1794 135
rect 1807 133 1812 135
rect 2054 132 2056 140
rect 1760 126 1765 128
rect 1779 127 1788 128
rect 1779 126 1783 127
rect 1782 123 1783 126
rect 1787 125 1788 127
rect 2050 131 2056 132
rect 2064 131 2066 140
rect 2074 131 2076 140
rect 2383 134 2385 142
rect 2050 127 2051 131
rect 2055 127 2056 131
rect 2070 130 2076 131
rect 2050 126 2056 127
rect 1787 123 1791 125
rect 1816 123 1821 125
rect 1782 122 1788 123
rect 1760 116 1765 118
rect 1779 116 1791 118
rect 1816 116 1821 118
rect 1474 103 1476 107
rect 583 90 585 95
rect 590 90 592 95
rect 1729 105 1735 106
rect 1729 103 1730 105
rect 1703 101 1708 103
rect 1718 101 1730 103
rect 1734 102 1735 105
rect 1782 108 1788 116
rect 1734 101 1738 102
rect 1729 100 1738 101
rect 1747 100 1752 102
rect 1782 104 1783 108
rect 1787 104 1788 108
rect 1697 96 1703 97
rect 1697 92 1698 96
rect 1702 93 1703 96
rect 1782 101 1788 104
rect 1782 98 1783 101
rect 1755 96 1759 98
rect 1779 97 1783 98
rect 1787 100 1788 101
rect 2054 113 2056 126
rect 2064 124 2066 127
rect 2070 126 2071 130
rect 2075 126 2076 130
rect 2379 133 2385 134
rect 2393 133 2395 142
rect 2403 133 2405 142
rect 2710 137 2712 145
rect 2379 129 2380 133
rect 2384 129 2385 133
rect 2399 132 2405 133
rect 2379 128 2385 129
rect 2070 125 2076 126
rect 2060 123 2066 124
rect 2060 119 2061 123
rect 2065 119 2066 123
rect 2060 118 2066 119
rect 2061 113 2063 118
rect 2074 116 2076 125
rect 1787 98 1791 100
rect 1819 98 1823 100
rect 1787 97 1788 98
rect 1779 96 1788 97
rect 1721 93 1738 95
rect 1747 93 1752 95
rect 1702 92 1708 93
rect 1697 91 1708 92
rect 1718 91 1724 93
rect 2383 115 2385 128
rect 2393 126 2395 129
rect 2399 128 2400 132
rect 2404 128 2405 132
rect 2706 136 2712 137
rect 2720 136 2722 145
rect 2730 136 2732 145
rect 2706 132 2707 136
rect 2711 132 2712 136
rect 2726 135 2732 136
rect 2706 131 2712 132
rect 2399 127 2405 128
rect 2389 125 2395 126
rect 2389 121 2390 125
rect 2394 121 2395 125
rect 2389 120 2395 121
rect 2390 115 2392 120
rect 2403 118 2405 127
rect 2710 118 2712 131
rect 2720 129 2722 132
rect 2726 131 2727 135
rect 2731 131 2732 135
rect 2726 130 2732 131
rect 2716 128 2722 129
rect 2716 124 2717 128
rect 2721 124 2722 128
rect 2716 123 2722 124
rect 2717 118 2719 123
rect 2730 121 2732 130
rect 2074 100 2076 104
rect 2403 102 2405 106
rect 2730 105 2732 109
rect 1782 91 1788 92
rect 1721 86 1727 87
rect 1721 83 1722 86
rect 1701 81 1706 83
rect 1718 82 1722 83
rect 1726 83 1727 86
rect 1755 89 1759 91
rect 1779 89 1783 91
rect 1782 87 1783 89
rect 1787 90 1788 91
rect 2054 91 2056 95
rect 2061 91 2063 95
rect 2383 93 2385 97
rect 2390 93 2392 97
rect 2710 96 2712 100
rect 2717 96 2719 100
rect 1787 88 1791 90
rect 1819 88 1827 90
rect 1787 87 1788 88
rect 1782 86 1788 87
rect 1726 82 1735 83
rect 1718 81 1735 82
rect 1741 81 1745 83
rect 1782 81 1788 82
rect 1782 80 1783 81
rect 1757 78 1759 80
rect 1773 78 1783 80
rect 1782 77 1783 78
rect 1787 80 1788 81
rect 1787 78 1791 80
rect 1819 78 1823 80
rect 1787 77 1788 78
rect 1782 76 1788 77
rect 1825 55 1827 88
rect 2255 68 2257 72
rect 2265 70 2267 75
rect 2275 70 2277 75
rect 1814 53 1827 55
rect 1814 16 1816 53
rect 2348 68 2350 72
rect 2358 70 2360 75
rect 2368 70 2370 75
rect 2255 46 2257 50
rect 2265 46 2267 57
rect 2275 54 2277 57
rect 2275 53 2281 54
rect 2275 49 2276 53
rect 2280 49 2281 53
rect 2435 68 2437 72
rect 2445 70 2447 75
rect 2455 70 2457 75
rect 2275 48 2281 49
rect 2255 45 2261 46
rect 2255 41 2256 45
rect 2260 41 2261 45
rect 2255 40 2261 41
rect 2265 45 2271 46
rect 2265 41 2266 45
rect 2270 41 2271 45
rect 2265 40 2271 41
rect 2255 35 2257 40
rect 2268 35 2270 40
rect 2275 35 2277 48
rect 2348 46 2350 50
rect 2358 46 2360 57
rect 2368 54 2370 57
rect 2368 53 2374 54
rect 2368 49 2369 53
rect 2373 49 2374 53
rect 2368 48 2374 49
rect 2348 45 2354 46
rect 2348 41 2349 45
rect 2353 41 2354 45
rect 2348 40 2354 41
rect 2358 45 2364 46
rect 2358 41 2359 45
rect 2363 41 2364 45
rect 2358 40 2364 41
rect 2348 35 2350 40
rect 2361 35 2363 40
rect 2368 35 2370 48
rect 2435 46 2437 50
rect 2445 46 2447 57
rect 2455 54 2457 57
rect 2455 53 2461 54
rect 2455 49 2456 53
rect 2460 49 2461 53
rect 2455 48 2461 49
rect 2435 45 2441 46
rect 2435 41 2436 45
rect 2440 41 2441 45
rect 2435 40 2441 41
rect 2445 45 2451 46
rect 2445 41 2446 45
rect 2450 41 2451 45
rect 2445 40 2451 41
rect 2435 35 2437 40
rect 2448 35 2450 40
rect 2455 35 2457 48
rect 2255 22 2257 26
rect 2268 19 2270 24
rect 2275 19 2277 24
rect 2348 22 2350 26
rect 2361 19 2363 24
rect 2368 19 2370 24
rect 2435 22 2437 26
rect 2448 19 2450 24
rect 2455 19 2457 24
<< ndiffusion >>
rect 1744 1056 1750 1057
rect 1744 1052 1745 1056
rect 1749 1055 1750 1056
rect 1749 1052 1753 1055
rect 1744 1050 1753 1052
rect 1744 1043 1753 1048
rect 1744 1039 1753 1041
rect 175 1029 182 1030
rect 175 1025 177 1029
rect 181 1025 182 1029
rect 175 1020 182 1025
rect 262 1029 269 1030
rect 262 1025 264 1029
rect 268 1025 269 1029
rect 157 1019 164 1020
rect 157 1015 158 1019
rect 162 1015 164 1019
rect 157 1014 164 1015
rect 159 1009 164 1014
rect 166 1009 171 1020
rect 173 1018 182 1020
rect 262 1020 269 1025
rect 355 1029 362 1030
rect 355 1025 357 1029
rect 361 1025 362 1029
rect 244 1019 251 1020
rect 173 1009 184 1018
rect 186 1017 193 1018
rect 186 1013 188 1017
rect 192 1013 193 1017
rect 244 1015 245 1019
rect 249 1015 251 1019
rect 244 1014 251 1015
rect 186 1012 193 1013
rect 186 1009 191 1012
rect 246 1009 251 1014
rect 253 1009 258 1020
rect 260 1018 269 1020
rect 355 1020 362 1025
rect 588 1031 595 1032
rect 588 1027 589 1031
rect 593 1027 595 1031
rect 337 1019 344 1020
rect 260 1009 271 1018
rect 273 1017 280 1018
rect 273 1013 275 1017
rect 279 1013 280 1017
rect 337 1015 338 1019
rect 342 1015 344 1019
rect 337 1014 344 1015
rect 273 1012 280 1013
rect 273 1009 278 1012
rect 339 1009 344 1014
rect 346 1009 351 1020
rect 353 1018 362 1020
rect 588 1022 595 1027
rect 681 1031 688 1032
rect 681 1027 682 1031
rect 686 1027 688 1031
rect 588 1020 597 1022
rect 577 1019 584 1020
rect 353 1009 364 1018
rect 366 1017 373 1018
rect 366 1013 368 1017
rect 372 1013 373 1017
rect 577 1015 578 1019
rect 582 1015 584 1019
rect 577 1014 584 1015
rect 366 1012 373 1013
rect 366 1009 371 1012
rect 579 1011 584 1014
rect 586 1011 597 1020
rect 599 1011 604 1022
rect 606 1021 613 1022
rect 606 1017 608 1021
rect 612 1017 613 1021
rect 681 1022 688 1027
rect 768 1031 775 1032
rect 768 1027 769 1031
rect 773 1027 775 1031
rect 1625 1028 1631 1029
rect 681 1020 690 1022
rect 606 1016 613 1017
rect 670 1019 677 1020
rect 606 1011 611 1016
rect 670 1015 671 1019
rect 675 1015 677 1019
rect 670 1014 677 1015
rect 672 1011 677 1014
rect 679 1011 690 1020
rect 692 1011 697 1022
rect 699 1021 706 1022
rect 699 1017 701 1021
rect 705 1017 706 1021
rect 768 1022 775 1027
rect 768 1020 777 1022
rect 699 1016 706 1017
rect 757 1019 764 1020
rect 699 1011 704 1016
rect 757 1015 758 1019
rect 762 1015 764 1019
rect 757 1014 764 1015
rect 759 1011 764 1014
rect 766 1011 777 1020
rect 779 1011 784 1022
rect 786 1021 793 1022
rect 786 1017 788 1021
rect 792 1017 793 1021
rect 786 1016 793 1017
rect 786 1011 791 1016
rect 1625 1024 1626 1028
rect 1630 1024 1631 1028
rect 1625 1022 1631 1024
rect 1741 1038 1759 1039
rect 1741 1034 1754 1038
rect 1758 1034 1759 1038
rect 1741 1033 1759 1034
rect 1741 1031 1747 1033
rect 1625 1018 1631 1020
rect 1613 1017 1631 1018
rect 1613 1013 1614 1017
rect 1618 1013 1631 1017
rect 1613 1012 1631 1013
rect 1741 1027 1747 1029
rect 1741 1023 1742 1027
rect 1746 1023 1747 1027
rect 1741 1022 1747 1023
rect 1619 1010 1628 1012
rect 1619 1003 1628 1008
rect 1619 999 1628 1001
rect 1619 996 1623 999
rect 1074 976 1085 979
rect 1087 976 1104 979
rect 1622 995 1623 996
rect 1627 995 1628 999
rect 1622 994 1628 995
rect 1741 1011 1759 1012
rect 1741 1007 1754 1011
rect 1758 1007 1759 1011
rect 1741 1006 1759 1007
rect 1741 1004 1753 1006
rect 1741 997 1753 1002
rect 1741 993 1753 995
rect 1741 989 1744 993
rect 1748 990 1753 993
rect 1748 989 1750 990
rect 1741 987 1750 989
rect 1186 980 1196 981
rect 1146 975 1157 978
rect 1159 975 1176 978
rect 1186 976 1188 980
rect 1192 976 1196 980
rect 1186 975 1196 976
rect 1198 975 1217 981
rect 1219 980 1227 981
rect 1219 976 1222 980
rect 1226 976 1227 980
rect 1219 975 1227 976
rect 1240 980 1250 981
rect 1240 976 1242 980
rect 1246 976 1250 980
rect 1240 975 1250 976
rect 1252 975 1271 981
rect 1273 980 1281 981
rect 1273 976 1276 980
rect 1280 976 1281 980
rect 1273 975 1281 976
rect 1296 980 1306 981
rect 1296 976 1298 980
rect 1302 976 1306 980
rect 1296 975 1306 976
rect 1308 975 1327 981
rect 1329 980 1337 981
rect 1329 976 1332 980
rect 1336 976 1337 980
rect 1329 975 1337 976
rect 1350 980 1360 981
rect 1350 976 1352 980
rect 1356 976 1360 980
rect 1350 975 1360 976
rect 1362 975 1381 981
rect 1383 980 1391 981
rect 1383 976 1386 980
rect 1390 976 1391 980
rect 1383 975 1391 976
rect 1741 983 1750 985
rect 1741 979 1742 983
rect 1746 979 1750 983
rect 1741 977 1750 979
rect 1741 971 1750 975
rect 1741 967 1745 971
rect 1749 967 1750 971
rect 1741 966 1750 967
rect 1736 961 1745 966
rect 79 902 86 903
rect 79 898 80 902
rect 84 898 86 902
rect 79 897 86 898
rect 88 900 96 903
rect 157 907 164 908
rect 157 903 158 907
rect 162 903 164 907
rect 157 902 164 903
rect 88 897 98 900
rect 90 891 98 897
rect 100 891 105 900
rect 107 899 114 900
rect 159 899 164 902
rect 166 903 171 908
rect 241 907 248 908
rect 241 903 242 907
rect 246 903 248 907
rect 166 899 180 903
rect 107 895 109 899
rect 113 895 114 899
rect 107 894 114 895
rect 171 895 172 899
rect 176 895 180 899
rect 171 894 180 895
rect 182 902 190 903
rect 182 898 184 902
rect 188 898 190 902
rect 182 894 190 898
rect 192 900 200 903
rect 192 896 194 900
rect 198 896 200 900
rect 192 894 200 896
rect 107 891 112 894
rect 90 890 96 891
rect 90 886 91 890
rect 95 886 96 890
rect 90 885 96 886
rect 195 891 200 894
rect 202 891 207 903
rect 209 891 217 903
rect 241 902 248 903
rect 243 899 248 902
rect 250 903 255 908
rect 250 899 264 903
rect 255 895 256 899
rect 260 895 264 899
rect 255 894 264 895
rect 266 902 274 903
rect 266 898 268 902
rect 272 898 274 902
rect 266 894 274 898
rect 276 900 284 903
rect 276 896 278 900
rect 282 896 284 900
rect 276 894 284 896
rect 211 890 217 891
rect 211 886 212 890
rect 216 886 217 890
rect 211 885 217 886
rect 279 891 284 894
rect 286 891 291 903
rect 293 891 301 903
rect 311 902 318 903
rect 311 898 312 902
rect 316 898 318 902
rect 311 897 318 898
rect 320 900 328 903
rect 408 904 415 905
rect 408 900 409 904
rect 413 900 415 904
rect 320 897 330 900
rect 322 891 330 897
rect 332 891 337 900
rect 339 899 346 900
rect 408 899 415 900
rect 417 902 425 905
rect 486 909 493 910
rect 486 905 487 909
rect 491 905 493 909
rect 486 904 493 905
rect 417 899 427 902
rect 339 895 341 899
rect 345 895 346 899
rect 339 894 346 895
rect 339 891 344 894
rect 419 893 427 899
rect 429 893 434 902
rect 436 901 443 902
rect 488 901 493 904
rect 495 905 500 910
rect 570 909 577 910
rect 570 905 571 909
rect 575 905 577 909
rect 495 901 509 905
rect 436 897 438 901
rect 442 897 443 901
rect 436 896 443 897
rect 500 897 501 901
rect 505 897 509 901
rect 500 896 509 897
rect 511 904 519 905
rect 511 900 513 904
rect 517 900 519 904
rect 511 896 519 900
rect 521 902 529 905
rect 521 898 523 902
rect 527 898 529 902
rect 521 896 529 898
rect 436 893 441 896
rect 295 890 301 891
rect 295 886 296 890
rect 300 886 301 890
rect 295 885 301 886
rect 322 890 328 891
rect 322 886 323 890
rect 327 886 328 890
rect 419 892 425 893
rect 419 888 420 892
rect 424 888 425 892
rect 419 887 425 888
rect 524 893 529 896
rect 531 893 536 905
rect 538 893 546 905
rect 570 904 577 905
rect 572 901 577 904
rect 579 905 584 910
rect 579 901 593 905
rect 584 897 585 901
rect 589 897 593 901
rect 584 896 593 897
rect 595 904 603 905
rect 595 900 597 904
rect 601 900 603 904
rect 595 896 603 900
rect 605 902 613 905
rect 605 898 607 902
rect 611 898 613 902
rect 605 896 613 898
rect 540 892 546 893
rect 540 888 541 892
rect 545 888 546 892
rect 540 887 546 888
rect 608 893 613 896
rect 615 893 620 905
rect 622 893 630 905
rect 640 904 647 905
rect 640 900 641 904
rect 645 900 647 904
rect 640 899 647 900
rect 649 902 657 905
rect 735 907 742 908
rect 735 903 736 907
rect 740 903 742 907
rect 735 902 742 903
rect 744 905 752 908
rect 1150 953 1161 956
rect 1163 953 1180 956
rect 1190 955 1200 956
rect 1190 951 1192 955
rect 1196 951 1200 955
rect 1190 950 1200 951
rect 1202 950 1221 956
rect 1223 955 1231 956
rect 1223 951 1226 955
rect 1230 951 1231 955
rect 1223 950 1231 951
rect 1244 955 1254 956
rect 1244 951 1246 955
rect 1250 951 1254 955
rect 1244 950 1254 951
rect 1256 950 1275 956
rect 1277 955 1285 956
rect 1277 951 1280 955
rect 1284 951 1285 955
rect 1277 950 1285 951
rect 1300 955 1310 956
rect 1300 951 1302 955
rect 1306 951 1310 955
rect 1300 950 1310 951
rect 1312 950 1331 956
rect 1333 955 1341 956
rect 1333 951 1336 955
rect 1340 951 1341 955
rect 1333 950 1341 951
rect 1354 955 1364 956
rect 1354 951 1356 955
rect 1360 951 1364 955
rect 1354 950 1364 951
rect 1366 950 1385 956
rect 1387 955 1395 956
rect 1387 951 1390 955
rect 1394 951 1395 955
rect 1736 957 1745 959
rect 1736 953 1737 957
rect 1741 954 1745 957
rect 1741 953 1742 954
rect 1736 952 1742 953
rect 1387 950 1395 951
rect 1630 950 1636 951
rect 1630 949 1631 950
rect 1627 946 1631 949
rect 1635 946 1636 950
rect 1627 944 1636 946
rect 813 912 820 913
rect 813 908 814 912
rect 818 908 820 912
rect 813 907 820 908
rect 744 902 754 905
rect 649 899 659 902
rect 651 893 659 899
rect 661 893 666 902
rect 668 901 675 902
rect 668 897 670 901
rect 674 897 675 901
rect 668 896 675 897
rect 746 896 754 902
rect 756 896 761 905
rect 763 904 770 905
rect 815 904 820 907
rect 822 908 827 913
rect 897 912 904 913
rect 897 908 898 912
rect 902 908 904 912
rect 822 904 836 908
rect 763 900 765 904
rect 769 900 770 904
rect 763 899 770 900
rect 827 900 828 904
rect 832 900 836 904
rect 827 899 836 900
rect 838 907 846 908
rect 838 903 840 907
rect 844 903 846 907
rect 838 899 846 903
rect 848 905 856 908
rect 848 901 850 905
rect 854 901 856 905
rect 848 899 856 901
rect 763 896 768 899
rect 668 893 673 896
rect 624 892 630 893
rect 624 888 625 892
rect 629 888 630 892
rect 624 887 630 888
rect 651 892 657 893
rect 651 888 652 892
rect 656 888 657 892
rect 746 895 752 896
rect 746 891 747 895
rect 751 891 752 895
rect 746 890 752 891
rect 851 896 856 899
rect 858 896 863 908
rect 865 896 873 908
rect 897 907 904 908
rect 899 904 904 907
rect 906 908 911 913
rect 906 904 920 908
rect 911 900 912 904
rect 916 900 920 904
rect 911 899 920 900
rect 922 907 930 908
rect 922 903 924 907
rect 928 903 930 907
rect 922 899 930 903
rect 932 905 940 908
rect 932 901 934 905
rect 938 901 940 905
rect 932 899 940 901
rect 867 895 873 896
rect 867 891 868 895
rect 872 891 873 895
rect 867 890 873 891
rect 935 896 940 899
rect 942 896 947 908
rect 949 896 957 908
rect 967 907 974 908
rect 967 903 968 907
rect 972 903 974 907
rect 967 902 974 903
rect 976 905 984 908
rect 1591 935 1597 936
rect 1591 931 1592 935
rect 1596 931 1597 935
rect 1591 929 1597 931
rect 1591 925 1597 927
rect 1591 921 1592 925
rect 1596 921 1597 925
rect 1591 919 1597 921
rect 1591 915 1597 917
rect 1591 911 1592 915
rect 1596 911 1597 915
rect 1591 909 1597 911
rect 976 902 986 905
rect 978 896 986 902
rect 988 896 993 905
rect 995 904 1002 905
rect 995 900 997 904
rect 1001 900 1002 904
rect 1591 905 1597 907
rect 1591 901 1592 905
rect 1596 901 1597 905
rect 1627 937 1636 942
rect 1622 936 1631 937
rect 1622 932 1623 936
rect 1627 932 1631 936
rect 1622 928 1631 932
rect 1622 924 1631 926
rect 1622 920 1626 924
rect 1630 920 1631 924
rect 1622 918 1631 920
rect 1741 927 1759 928
rect 1741 923 1754 927
rect 1758 923 1759 927
rect 1741 922 1759 923
rect 1741 920 1753 922
rect 1622 914 1631 916
rect 1622 913 1624 914
rect 1619 910 1624 913
rect 1628 910 1631 914
rect 1619 908 1631 910
rect 1775 918 1781 919
rect 1741 913 1753 918
rect 1619 901 1631 906
rect 1591 900 1597 901
rect 995 899 1002 900
rect 1741 909 1753 911
rect 1741 905 1744 909
rect 1748 906 1753 909
rect 1748 905 1750 906
rect 1741 903 1750 905
rect 995 896 1000 899
rect 1619 897 1631 899
rect 1613 896 1631 897
rect 951 895 957 896
rect 951 891 952 895
rect 956 891 957 895
rect 951 890 957 891
rect 978 895 984 896
rect 978 891 979 895
rect 983 891 984 895
rect 1613 892 1614 896
rect 1618 892 1631 896
rect 978 890 984 891
rect 651 887 657 888
rect 322 885 328 886
rect 1613 891 1631 892
rect 1741 899 1750 901
rect 1741 895 1742 899
rect 1746 895 1750 899
rect 1741 893 1750 895
rect 828 873 835 874
rect 501 870 508 871
rect 172 868 179 869
rect 172 864 173 868
rect 177 864 179 868
rect 172 863 179 864
rect 181 868 189 869
rect 181 864 183 868
rect 187 864 189 868
rect 181 863 189 864
rect 191 868 199 869
rect 191 864 193 868
rect 197 864 199 868
rect 191 863 199 864
rect 201 868 208 869
rect 201 864 203 868
rect 207 864 208 868
rect 501 866 502 870
rect 506 866 508 870
rect 501 865 508 866
rect 510 870 518 871
rect 510 866 512 870
rect 516 866 518 870
rect 510 865 518 866
rect 520 870 528 871
rect 520 866 522 870
rect 526 866 528 870
rect 520 865 528 866
rect 530 870 537 871
rect 530 866 532 870
rect 536 866 537 870
rect 828 869 829 873
rect 833 869 835 873
rect 828 868 835 869
rect 837 873 845 874
rect 837 869 839 873
rect 843 869 845 873
rect 837 868 845 869
rect 847 873 855 874
rect 847 869 849 873
rect 853 869 855 873
rect 847 868 855 869
rect 857 873 864 874
rect 857 869 859 873
rect 863 869 864 873
rect 857 868 864 869
rect 530 865 537 866
rect 201 863 208 864
rect 1741 887 1750 891
rect 1741 883 1745 887
rect 1749 883 1750 887
rect 1741 882 1750 883
rect 1736 877 1745 882
rect 1775 914 1776 918
rect 1780 914 1781 918
rect 1775 912 1781 914
rect 1775 908 1781 910
rect 1775 904 1776 908
rect 1780 904 1781 908
rect 1775 902 1781 904
rect 1775 898 1781 900
rect 1775 894 1776 898
rect 1780 894 1781 898
rect 1775 892 1781 894
rect 1775 888 1781 890
rect 1775 884 1776 888
rect 1780 884 1781 888
rect 1775 883 1781 884
rect 2700 883 2705 890
rect 2451 882 2458 883
rect 2451 878 2452 882
rect 2456 878 2458 882
rect 2451 877 2458 878
rect 2460 882 2468 883
rect 2460 878 2462 882
rect 2466 878 2468 882
rect 2460 877 2468 878
rect 2470 882 2478 883
rect 2470 878 2472 882
rect 2476 878 2478 882
rect 2470 877 2478 878
rect 2480 882 2487 883
rect 2480 878 2482 882
rect 2486 878 2487 882
rect 2480 877 2487 878
rect 2678 882 2685 883
rect 2678 878 2679 882
rect 2683 878 2685 882
rect 2678 877 2685 878
rect 1736 873 1745 875
rect 1736 869 1737 873
rect 1741 870 1745 873
rect 1741 869 1742 870
rect 2680 870 2685 877
rect 2687 878 2695 883
rect 2687 874 2689 878
rect 2693 874 2695 878
rect 2687 873 2695 874
rect 2697 881 2705 883
rect 2697 877 2699 881
rect 2703 877 2705 881
rect 2697 876 2705 877
rect 2707 889 2715 890
rect 2707 885 2709 889
rect 2713 885 2715 889
rect 2707 876 2715 885
rect 2717 889 2724 890
rect 2717 885 2719 889
rect 2723 885 2724 889
rect 2717 882 2724 885
rect 2730 883 2735 890
rect 2717 878 2719 882
rect 2723 878 2724 882
rect 2717 876 2724 878
rect 2728 882 2735 883
rect 2728 878 2729 882
rect 2733 878 2735 882
rect 2728 877 2735 878
rect 2697 873 2702 876
rect 2687 870 2692 873
rect 1736 868 1742 869
rect 1630 866 1636 867
rect 1630 865 1631 866
rect 1627 862 1631 865
rect 1635 862 1636 866
rect 1627 860 1636 862
rect 2730 870 2735 877
rect 2737 870 2742 890
rect 2744 884 2751 890
rect 2811 884 2818 885
rect 2744 875 2753 884
rect 2744 871 2746 875
rect 2750 871 2753 875
rect 2744 870 2753 871
rect 2755 882 2762 884
rect 2755 878 2757 882
rect 2761 878 2762 882
rect 2811 880 2812 884
rect 2816 880 2818 884
rect 2811 879 2818 880
rect 2820 884 2828 885
rect 2820 880 2822 884
rect 2826 880 2828 884
rect 2820 879 2828 880
rect 2830 884 2838 885
rect 2830 880 2832 884
rect 2836 880 2838 884
rect 2830 879 2838 880
rect 2840 884 2847 885
rect 2840 880 2842 884
rect 2846 880 2847 884
rect 2840 879 2847 880
rect 2755 877 2762 878
rect 2755 870 2760 877
rect 2691 862 2697 863
rect 2331 860 2337 861
rect 1074 831 1085 834
rect 1087 831 1104 834
rect 1419 847 1426 848
rect 1419 843 1420 847
rect 1424 843 1426 847
rect 1419 842 1426 843
rect 1421 838 1426 842
rect 1428 839 1438 848
rect 1428 838 1431 839
rect 1186 835 1196 836
rect 1146 830 1157 833
rect 1159 830 1176 833
rect 1186 831 1188 835
rect 1192 831 1196 835
rect 1186 830 1196 831
rect 1198 830 1217 836
rect 1219 835 1227 836
rect 1219 831 1222 835
rect 1226 831 1227 835
rect 1219 830 1227 831
rect 1240 835 1250 836
rect 1240 831 1242 835
rect 1246 831 1250 835
rect 1240 830 1250 831
rect 1252 830 1271 836
rect 1273 835 1281 836
rect 1273 831 1276 835
rect 1280 831 1281 835
rect 1273 830 1281 831
rect 1296 835 1306 836
rect 1296 831 1298 835
rect 1302 831 1306 835
rect 1296 830 1306 831
rect 1308 830 1327 836
rect 1329 835 1337 836
rect 1329 831 1332 835
rect 1336 831 1337 835
rect 1329 830 1337 831
rect 1350 835 1360 836
rect 1350 831 1352 835
rect 1356 831 1360 835
rect 1350 830 1360 831
rect 1362 830 1381 836
rect 1383 835 1391 836
rect 1383 831 1386 835
rect 1390 831 1391 835
rect 1430 835 1431 838
rect 1435 835 1438 839
rect 1430 834 1438 835
rect 1440 847 1447 848
rect 1440 843 1442 847
rect 1446 843 1447 847
rect 1440 840 1447 843
rect 1440 836 1442 840
rect 1446 836 1447 840
rect 1440 834 1447 836
rect 1627 853 1636 858
rect 1622 852 1631 853
rect 1622 848 1623 852
rect 1627 848 1631 852
rect 2331 856 2332 860
rect 2336 856 2337 860
rect 2331 855 2337 856
rect 2358 860 2364 861
rect 2358 856 2359 860
rect 2363 856 2364 860
rect 2358 855 2364 856
rect 2315 852 2320 855
rect 1622 844 1631 848
rect 2313 851 2320 852
rect 2313 847 2314 851
rect 2318 847 2320 851
rect 2313 846 2320 847
rect 2322 846 2327 855
rect 2329 849 2337 855
rect 2329 846 2339 849
rect 1622 840 1631 842
rect 1622 836 1626 840
rect 1630 836 1631 840
rect 1622 834 1631 836
rect 1383 830 1391 831
rect 1622 830 1631 832
rect 1622 829 1624 830
rect 1619 826 1624 829
rect 1628 826 1631 830
rect 1619 824 1631 826
rect 2331 843 2339 846
rect 2341 848 2348 849
rect 2341 844 2343 848
rect 2347 844 2348 848
rect 2341 843 2348 844
rect 2358 843 2366 855
rect 2368 843 2373 855
rect 2375 852 2380 855
rect 2442 860 2448 861
rect 2442 856 2443 860
rect 2447 856 2448 860
rect 2442 855 2448 856
rect 2375 850 2383 852
rect 2375 846 2377 850
rect 2381 846 2383 850
rect 2375 843 2383 846
rect 2385 848 2393 852
rect 2385 844 2387 848
rect 2391 844 2393 848
rect 2385 843 2393 844
rect 2395 851 2404 852
rect 2395 847 2399 851
rect 2403 847 2404 851
rect 2395 843 2409 847
rect 2404 838 2409 843
rect 2411 844 2416 847
rect 2411 843 2418 844
rect 2442 843 2450 855
rect 2452 843 2457 855
rect 2459 852 2464 855
rect 2563 860 2569 861
rect 2563 856 2564 860
rect 2568 856 2569 860
rect 2563 855 2569 856
rect 2691 858 2692 862
rect 2696 858 2697 862
rect 2691 857 2697 858
rect 2718 862 2724 863
rect 2718 858 2719 862
rect 2723 858 2724 862
rect 2718 857 2724 858
rect 2547 852 2552 855
rect 2459 850 2467 852
rect 2459 846 2461 850
rect 2465 846 2467 850
rect 2459 843 2467 846
rect 2469 848 2477 852
rect 2469 844 2471 848
rect 2475 844 2477 848
rect 2469 843 2477 844
rect 2479 851 2488 852
rect 2479 847 2483 851
rect 2487 847 2488 851
rect 2545 851 2552 852
rect 2545 847 2546 851
rect 2550 847 2552 851
rect 2479 843 2493 847
rect 2411 839 2413 843
rect 2417 839 2418 843
rect 2411 838 2418 839
rect 2488 838 2493 843
rect 2495 844 2500 847
rect 2545 846 2552 847
rect 2554 846 2559 855
rect 2561 849 2569 855
rect 2675 854 2680 857
rect 2673 853 2680 854
rect 2673 849 2674 853
rect 2678 849 2680 853
rect 2561 846 2571 849
rect 2495 843 2502 844
rect 2495 839 2497 843
rect 2501 839 2502 843
rect 2495 838 2502 839
rect 78 756 85 757
rect 78 752 79 756
rect 83 752 85 756
rect 78 751 85 752
rect 87 754 95 757
rect 156 761 163 762
rect 156 757 157 761
rect 161 757 163 761
rect 156 756 163 757
rect 87 751 97 754
rect 89 745 97 751
rect 99 745 104 754
rect 106 753 113 754
rect 158 753 163 756
rect 165 757 170 762
rect 240 761 247 762
rect 240 757 241 761
rect 245 757 247 761
rect 165 753 179 757
rect 106 749 108 753
rect 112 749 113 753
rect 106 748 113 749
rect 170 749 171 753
rect 175 749 179 753
rect 170 748 179 749
rect 181 756 189 757
rect 181 752 183 756
rect 187 752 189 756
rect 181 748 189 752
rect 191 754 199 757
rect 191 750 193 754
rect 197 750 199 754
rect 191 748 199 750
rect 106 745 111 748
rect 89 744 95 745
rect 89 740 90 744
rect 94 740 95 744
rect 89 739 95 740
rect 194 745 199 748
rect 201 745 206 757
rect 208 745 216 757
rect 240 756 247 757
rect 242 753 247 756
rect 249 757 254 762
rect 249 753 263 757
rect 254 749 255 753
rect 259 749 263 753
rect 254 748 263 749
rect 265 756 273 757
rect 265 752 267 756
rect 271 752 273 756
rect 265 748 273 752
rect 275 754 283 757
rect 275 750 277 754
rect 281 750 283 754
rect 275 748 283 750
rect 210 744 216 745
rect 210 740 211 744
rect 215 740 216 744
rect 210 739 216 740
rect 278 745 283 748
rect 285 745 290 757
rect 292 745 300 757
rect 310 756 317 757
rect 310 752 311 756
rect 315 752 317 756
rect 310 751 317 752
rect 319 754 327 757
rect 407 758 414 759
rect 407 754 408 758
rect 412 754 414 758
rect 319 751 329 754
rect 321 745 329 751
rect 331 745 336 754
rect 338 753 345 754
rect 407 753 414 754
rect 416 756 424 759
rect 485 763 492 764
rect 485 759 486 763
rect 490 759 492 763
rect 485 758 492 759
rect 416 753 426 756
rect 338 749 340 753
rect 344 749 345 753
rect 338 748 345 749
rect 338 745 343 748
rect 418 747 426 753
rect 428 747 433 756
rect 435 755 442 756
rect 487 755 492 758
rect 494 759 499 764
rect 569 763 576 764
rect 569 759 570 763
rect 574 759 576 763
rect 494 755 508 759
rect 435 751 437 755
rect 441 751 442 755
rect 435 750 442 751
rect 499 751 500 755
rect 504 751 508 755
rect 499 750 508 751
rect 510 758 518 759
rect 510 754 512 758
rect 516 754 518 758
rect 510 750 518 754
rect 520 756 528 759
rect 520 752 522 756
rect 526 752 528 756
rect 520 750 528 752
rect 435 747 440 750
rect 294 744 300 745
rect 294 740 295 744
rect 299 740 300 744
rect 294 739 300 740
rect 321 744 327 745
rect 321 740 322 744
rect 326 740 327 744
rect 418 746 424 747
rect 418 742 419 746
rect 423 742 424 746
rect 418 741 424 742
rect 523 747 528 750
rect 530 747 535 759
rect 537 747 545 759
rect 569 758 576 759
rect 571 755 576 758
rect 578 759 583 764
rect 578 755 592 759
rect 583 751 584 755
rect 588 751 592 755
rect 583 750 592 751
rect 594 758 602 759
rect 594 754 596 758
rect 600 754 602 758
rect 594 750 602 754
rect 604 756 612 759
rect 604 752 606 756
rect 610 752 612 756
rect 604 750 612 752
rect 539 746 545 747
rect 539 742 540 746
rect 544 742 545 746
rect 539 741 545 742
rect 607 747 612 750
rect 614 747 619 759
rect 621 747 629 759
rect 639 758 646 759
rect 639 754 640 758
rect 644 754 646 758
rect 639 753 646 754
rect 648 756 656 759
rect 734 761 741 762
rect 734 757 735 761
rect 739 757 741 761
rect 734 756 741 757
rect 743 759 751 762
rect 1150 808 1161 811
rect 1163 808 1180 811
rect 1190 810 1200 811
rect 1190 806 1192 810
rect 1196 806 1200 810
rect 1190 805 1200 806
rect 1202 805 1221 811
rect 1223 810 1231 811
rect 1223 806 1226 810
rect 1230 806 1231 810
rect 1223 805 1231 806
rect 1244 810 1254 811
rect 1244 806 1246 810
rect 1250 806 1254 810
rect 1244 805 1254 806
rect 1256 805 1275 811
rect 1277 810 1285 811
rect 1277 806 1280 810
rect 1284 806 1285 810
rect 1277 805 1285 806
rect 1300 810 1310 811
rect 1300 806 1302 810
rect 1306 806 1310 810
rect 1300 805 1310 806
rect 1312 805 1331 811
rect 1333 810 1341 811
rect 1333 806 1336 810
rect 1340 806 1341 810
rect 1333 805 1341 806
rect 1354 810 1364 811
rect 1354 806 1356 810
rect 1360 806 1364 810
rect 1354 805 1364 806
rect 1366 805 1385 811
rect 1387 810 1395 811
rect 1387 806 1390 810
rect 1394 806 1395 810
rect 1619 817 1631 822
rect 1619 813 1631 815
rect 1431 812 1439 813
rect 1431 809 1432 812
rect 1387 805 1395 806
rect 1422 805 1427 809
rect 1420 804 1427 805
rect 1420 800 1421 804
rect 1425 800 1427 804
rect 1420 799 1427 800
rect 1429 808 1432 809
rect 1436 808 1439 812
rect 1429 799 1439 808
rect 1441 811 1448 813
rect 1441 807 1443 811
rect 1447 807 1448 811
rect 1613 812 1631 813
rect 1613 808 1614 812
rect 1618 808 1631 812
rect 1613 807 1631 808
rect 1744 824 1750 825
rect 1744 820 1745 824
rect 1749 823 1750 824
rect 1749 820 1753 823
rect 1744 818 1753 820
rect 1441 804 1448 807
rect 1441 800 1443 804
rect 1447 800 1448 804
rect 1441 799 1448 800
rect 1744 811 1753 816
rect 1744 807 1753 809
rect 1625 796 1631 797
rect 1625 792 1626 796
rect 1630 792 1631 796
rect 1625 790 1631 792
rect 1741 806 1759 807
rect 1741 802 1754 806
rect 1758 802 1759 806
rect 1741 801 1759 802
rect 1741 799 1747 801
rect 812 766 819 767
rect 812 762 813 766
rect 817 762 819 766
rect 812 761 819 762
rect 743 756 753 759
rect 648 753 658 756
rect 650 747 658 753
rect 660 747 665 756
rect 667 755 674 756
rect 667 751 669 755
rect 673 751 674 755
rect 667 750 674 751
rect 745 750 753 756
rect 755 750 760 759
rect 762 758 769 759
rect 814 758 819 761
rect 821 762 826 767
rect 896 766 903 767
rect 896 762 897 766
rect 901 762 903 766
rect 821 758 835 762
rect 762 754 764 758
rect 768 754 769 758
rect 762 753 769 754
rect 826 754 827 758
rect 831 754 835 758
rect 826 753 835 754
rect 837 761 845 762
rect 837 757 839 761
rect 843 757 845 761
rect 837 753 845 757
rect 847 759 855 762
rect 847 755 849 759
rect 853 755 855 759
rect 847 753 855 755
rect 762 750 767 753
rect 667 747 672 750
rect 623 746 629 747
rect 623 742 624 746
rect 628 742 629 746
rect 623 741 629 742
rect 650 746 656 747
rect 650 742 651 746
rect 655 742 656 746
rect 745 749 751 750
rect 745 745 746 749
rect 750 745 751 749
rect 745 744 751 745
rect 850 750 855 753
rect 857 750 862 762
rect 864 750 872 762
rect 896 761 903 762
rect 898 758 903 761
rect 905 762 910 767
rect 905 758 919 762
rect 910 754 911 758
rect 915 754 919 758
rect 910 753 919 754
rect 921 761 929 762
rect 921 757 923 761
rect 927 757 929 761
rect 921 753 929 757
rect 931 759 939 762
rect 931 755 933 759
rect 937 755 939 759
rect 931 753 939 755
rect 866 749 872 750
rect 866 745 867 749
rect 871 745 872 749
rect 866 744 872 745
rect 934 750 939 753
rect 941 750 946 762
rect 948 750 956 762
rect 966 761 973 762
rect 966 757 967 761
rect 971 757 973 761
rect 966 756 973 757
rect 975 759 983 762
rect 975 756 985 759
rect 977 750 985 756
rect 987 750 992 759
rect 994 758 1001 759
rect 994 754 996 758
rect 1000 754 1001 758
rect 1625 786 1631 788
rect 1613 785 1631 786
rect 1613 781 1614 785
rect 1618 781 1631 785
rect 1613 780 1631 781
rect 1741 795 1747 797
rect 1741 791 1742 795
rect 1746 791 1747 795
rect 2563 843 2571 846
rect 2573 848 2580 849
rect 2673 848 2680 849
rect 2682 848 2687 857
rect 2689 851 2697 857
rect 2689 848 2699 851
rect 2573 844 2575 848
rect 2579 844 2580 848
rect 2573 843 2580 844
rect 2691 845 2699 848
rect 2701 850 2708 851
rect 2701 846 2703 850
rect 2707 846 2708 850
rect 2701 845 2708 846
rect 2718 845 2726 857
rect 2728 845 2733 857
rect 2735 854 2740 857
rect 2802 862 2808 863
rect 2802 858 2803 862
rect 2807 858 2808 862
rect 2802 857 2808 858
rect 2735 852 2743 854
rect 2735 848 2737 852
rect 2741 848 2743 852
rect 2735 845 2743 848
rect 2745 850 2753 854
rect 2745 846 2747 850
rect 2751 846 2753 850
rect 2745 845 2753 846
rect 2755 853 2764 854
rect 2755 849 2759 853
rect 2763 849 2764 853
rect 2755 845 2769 849
rect 2764 840 2769 845
rect 2771 846 2776 849
rect 2771 845 2778 846
rect 2802 845 2810 857
rect 2812 845 2817 857
rect 2819 854 2824 857
rect 2923 862 2929 863
rect 2923 858 2924 862
rect 2928 858 2929 862
rect 2923 857 2929 858
rect 2907 854 2912 857
rect 2819 852 2827 854
rect 2819 848 2821 852
rect 2825 848 2827 852
rect 2819 845 2827 848
rect 2829 850 2837 854
rect 2829 846 2831 850
rect 2835 846 2837 850
rect 2829 845 2837 846
rect 2839 853 2848 854
rect 2839 849 2843 853
rect 2847 849 2848 853
rect 2905 853 2912 854
rect 2905 849 2906 853
rect 2910 849 2912 853
rect 2839 845 2853 849
rect 2771 841 2773 845
rect 2777 841 2778 845
rect 2771 840 2778 841
rect 2848 840 2853 845
rect 2855 846 2860 849
rect 2905 848 2912 849
rect 2914 848 2919 857
rect 2921 851 2929 857
rect 2921 848 2931 851
rect 2855 845 2862 846
rect 2855 841 2857 845
rect 2861 841 2862 845
rect 2855 840 2862 841
rect 2923 845 2931 848
rect 2933 850 2940 851
rect 2933 846 2935 850
rect 2939 846 2940 850
rect 2933 845 2940 846
rect 1741 790 1747 791
rect 1619 778 1628 780
rect 1619 771 1628 776
rect 1619 767 1628 769
rect 1619 764 1623 767
rect 1622 763 1623 764
rect 1627 763 1628 767
rect 1622 762 1628 763
rect 994 753 1001 754
rect 994 750 999 753
rect 950 749 956 750
rect 950 745 951 749
rect 955 745 956 749
rect 950 744 956 745
rect 977 749 983 750
rect 977 745 978 749
rect 982 745 983 749
rect 977 744 983 745
rect 650 741 656 742
rect 321 739 327 740
rect 827 727 834 728
rect 500 724 507 725
rect 171 722 178 723
rect 171 718 172 722
rect 176 718 178 722
rect 171 717 178 718
rect 180 722 188 723
rect 180 718 182 722
rect 186 718 188 722
rect 180 717 188 718
rect 190 722 198 723
rect 190 718 192 722
rect 196 718 198 722
rect 190 717 198 718
rect 200 722 207 723
rect 200 718 202 722
rect 206 718 207 722
rect 500 720 501 724
rect 505 720 507 724
rect 500 719 507 720
rect 509 724 517 725
rect 509 720 511 724
rect 515 720 517 724
rect 509 719 517 720
rect 519 724 527 725
rect 519 720 521 724
rect 525 720 527 724
rect 519 719 527 720
rect 529 724 536 725
rect 529 720 531 724
rect 535 720 536 724
rect 827 723 828 727
rect 832 723 834 727
rect 827 722 834 723
rect 836 727 844 728
rect 836 723 838 727
rect 842 723 844 727
rect 836 722 844 723
rect 846 727 854 728
rect 846 723 848 727
rect 852 723 854 727
rect 846 722 854 723
rect 856 727 863 728
rect 856 723 858 727
rect 862 723 863 727
rect 856 722 863 723
rect 529 719 536 720
rect 200 717 207 718
rect 1985 740 1992 741
rect 1985 736 1986 740
rect 1990 736 1992 740
rect 1985 735 1992 736
rect 1994 738 2002 741
rect 2063 745 2070 746
rect 2063 741 2064 745
rect 2068 741 2070 745
rect 2063 740 2070 741
rect 1994 735 2004 738
rect 1996 729 2004 735
rect 2006 729 2011 738
rect 2013 737 2020 738
rect 2065 737 2070 740
rect 2072 741 2077 746
rect 2147 745 2154 746
rect 2147 741 2148 745
rect 2152 741 2154 745
rect 2072 737 2086 741
rect 2013 733 2015 737
rect 2019 733 2020 737
rect 2013 732 2020 733
rect 2077 733 2078 737
rect 2082 733 2086 737
rect 2077 732 2086 733
rect 2088 740 2096 741
rect 2088 736 2090 740
rect 2094 736 2096 740
rect 2088 732 2096 736
rect 2098 738 2106 741
rect 2098 734 2100 738
rect 2104 734 2106 738
rect 2098 732 2106 734
rect 2013 729 2018 732
rect 1996 728 2002 729
rect 1996 724 1997 728
rect 2001 724 2002 728
rect 1996 723 2002 724
rect 2101 729 2106 732
rect 2108 729 2113 741
rect 2115 729 2123 741
rect 2147 740 2154 741
rect 2149 737 2154 740
rect 2156 741 2161 746
rect 2156 737 2170 741
rect 2161 733 2162 737
rect 2166 733 2170 737
rect 2161 732 2170 733
rect 2172 740 2180 741
rect 2172 736 2174 740
rect 2178 736 2180 740
rect 2172 732 2180 736
rect 2182 738 2190 741
rect 2182 734 2184 738
rect 2188 734 2190 738
rect 2182 732 2190 734
rect 2117 728 2123 729
rect 2117 724 2118 728
rect 2122 724 2123 728
rect 2117 723 2123 724
rect 2185 729 2190 732
rect 2192 729 2197 741
rect 2199 729 2207 741
rect 2217 740 2224 741
rect 2217 736 2218 740
rect 2222 736 2224 740
rect 2217 735 2224 736
rect 2226 738 2234 741
rect 2226 735 2236 738
rect 2228 729 2236 735
rect 2238 729 2243 738
rect 2245 737 2252 738
rect 2245 733 2247 737
rect 2251 733 2252 737
rect 2245 732 2252 733
rect 2341 732 2348 733
rect 2245 729 2250 732
rect 2201 728 2207 729
rect 2201 724 2202 728
rect 2206 724 2207 728
rect 2201 723 2207 724
rect 2228 728 2234 729
rect 2228 724 2229 728
rect 2233 724 2234 728
rect 2341 728 2342 732
rect 2346 728 2348 732
rect 2341 727 2348 728
rect 2350 730 2358 733
rect 2419 737 2426 738
rect 2419 733 2420 737
rect 2424 733 2426 737
rect 2419 732 2426 733
rect 2350 727 2360 730
rect 2228 723 2234 724
rect 2352 721 2360 727
rect 2362 721 2367 730
rect 2369 729 2376 730
rect 2421 729 2426 732
rect 2428 733 2433 738
rect 2503 737 2510 738
rect 2503 733 2504 737
rect 2508 733 2510 737
rect 2428 729 2442 733
rect 2369 725 2371 729
rect 2375 725 2376 729
rect 2369 724 2376 725
rect 2433 725 2434 729
rect 2438 725 2442 729
rect 2433 724 2442 725
rect 2444 732 2452 733
rect 2444 728 2446 732
rect 2450 728 2452 732
rect 2444 724 2452 728
rect 2454 730 2462 733
rect 2454 726 2456 730
rect 2460 726 2462 730
rect 2454 724 2462 726
rect 2369 721 2374 724
rect 1073 689 1084 692
rect 1086 689 1103 692
rect 1984 710 1989 717
rect 1982 709 1989 710
rect 1419 707 1426 708
rect 1419 703 1420 707
rect 1424 703 1426 707
rect 1419 702 1426 703
rect 1421 698 1426 702
rect 1428 699 1438 708
rect 1428 698 1431 699
rect 1185 693 1195 694
rect 1145 688 1156 691
rect 1158 688 1175 691
rect 1185 689 1187 693
rect 1191 689 1195 693
rect 1185 688 1195 689
rect 1197 688 1216 694
rect 1218 693 1226 694
rect 1218 689 1221 693
rect 1225 689 1226 693
rect 1218 688 1226 689
rect 1239 693 1249 694
rect 1239 689 1241 693
rect 1245 689 1249 693
rect 1239 688 1249 689
rect 1251 688 1270 694
rect 1272 693 1280 694
rect 1272 689 1275 693
rect 1279 689 1280 693
rect 1272 688 1280 689
rect 1295 693 1305 694
rect 1295 689 1297 693
rect 1301 689 1305 693
rect 1295 688 1305 689
rect 1307 688 1326 694
rect 1328 693 1336 694
rect 1328 689 1331 693
rect 1335 689 1336 693
rect 1328 688 1336 689
rect 1349 693 1359 694
rect 1349 689 1351 693
rect 1355 689 1359 693
rect 1349 688 1359 689
rect 1361 688 1380 694
rect 1382 693 1390 694
rect 1430 695 1431 698
rect 1435 695 1438 699
rect 1430 694 1438 695
rect 1440 707 1447 708
rect 1440 703 1442 707
rect 1446 703 1447 707
rect 1982 705 1983 709
rect 1987 705 1989 709
rect 1982 703 1989 705
rect 1991 716 2000 717
rect 1991 712 1994 716
rect 1998 712 2000 716
rect 1991 703 2000 712
rect 1440 700 1447 703
rect 1440 696 1442 700
rect 1446 696 1447 700
rect 1440 694 1447 696
rect 1382 689 1385 693
rect 1389 689 1390 693
rect 1382 688 1390 689
rect 1746 696 1752 697
rect 1746 692 1747 696
rect 1751 695 1752 696
rect 1751 692 1755 695
rect 1993 697 2000 703
rect 2002 697 2007 717
rect 2009 710 2014 717
rect 2052 714 2057 717
rect 2042 711 2047 714
rect 2009 709 2016 710
rect 2009 705 2011 709
rect 2015 705 2016 709
rect 2009 704 2016 705
rect 2020 709 2027 711
rect 2020 705 2021 709
rect 2025 705 2027 709
rect 2009 697 2014 704
rect 2020 702 2027 705
rect 2020 698 2021 702
rect 2025 698 2027 702
rect 2020 697 2027 698
rect 2029 702 2037 711
rect 2029 698 2031 702
rect 2035 698 2037 702
rect 2029 697 2037 698
rect 2039 710 2047 711
rect 2039 706 2041 710
rect 2045 706 2047 710
rect 2039 704 2047 706
rect 2049 713 2057 714
rect 2049 709 2051 713
rect 2055 709 2057 713
rect 2049 704 2057 709
rect 2059 710 2064 717
rect 2352 720 2358 721
rect 2352 716 2353 720
rect 2357 716 2358 720
rect 2352 715 2358 716
rect 2457 721 2462 724
rect 2464 721 2469 733
rect 2471 721 2479 733
rect 2503 732 2510 733
rect 2505 729 2510 732
rect 2512 733 2517 738
rect 2512 729 2526 733
rect 2517 725 2518 729
rect 2522 725 2526 729
rect 2517 724 2526 725
rect 2528 732 2536 733
rect 2528 728 2530 732
rect 2534 728 2536 732
rect 2528 724 2536 728
rect 2538 730 2546 733
rect 2538 726 2540 730
rect 2544 726 2546 730
rect 2538 724 2546 726
rect 2473 720 2479 721
rect 2473 716 2474 720
rect 2478 716 2479 720
rect 2473 715 2479 716
rect 2541 721 2546 724
rect 2548 721 2553 733
rect 2555 721 2563 733
rect 2573 732 2580 733
rect 2573 728 2574 732
rect 2578 728 2580 732
rect 2573 727 2580 728
rect 2582 730 2590 733
rect 2701 734 2708 735
rect 2701 730 2702 734
rect 2706 730 2708 734
rect 2582 727 2592 730
rect 2584 721 2592 727
rect 2594 721 2599 730
rect 2601 729 2608 730
rect 2701 729 2708 730
rect 2710 732 2718 735
rect 2779 739 2786 740
rect 2779 735 2780 739
rect 2784 735 2786 739
rect 2779 734 2786 735
rect 2710 729 2720 732
rect 2601 725 2603 729
rect 2607 725 2608 729
rect 2601 724 2608 725
rect 2601 721 2606 724
rect 2712 723 2720 729
rect 2722 723 2727 732
rect 2729 731 2736 732
rect 2781 731 2786 734
rect 2788 735 2793 740
rect 2863 739 2870 740
rect 2863 735 2864 739
rect 2868 735 2870 739
rect 2788 731 2802 735
rect 2729 727 2731 731
rect 2735 727 2736 731
rect 2729 726 2736 727
rect 2793 727 2794 731
rect 2798 727 2802 731
rect 2793 726 2802 727
rect 2804 734 2812 735
rect 2804 730 2806 734
rect 2810 730 2812 734
rect 2804 726 2812 730
rect 2814 732 2822 735
rect 2814 728 2816 732
rect 2820 728 2822 732
rect 2814 726 2822 728
rect 2729 723 2734 726
rect 2557 720 2563 721
rect 2557 716 2558 720
rect 2562 716 2563 720
rect 2557 715 2563 716
rect 2584 720 2590 721
rect 2584 716 2585 720
rect 2589 716 2590 720
rect 2712 722 2718 723
rect 2712 718 2713 722
rect 2717 718 2718 722
rect 2712 717 2718 718
rect 2817 723 2822 726
rect 2824 723 2829 735
rect 2831 723 2839 735
rect 2863 734 2870 735
rect 2865 731 2870 734
rect 2872 735 2877 740
rect 2872 731 2886 735
rect 2877 727 2878 731
rect 2882 727 2886 731
rect 2877 726 2886 727
rect 2888 734 2896 735
rect 2888 730 2890 734
rect 2894 730 2896 734
rect 2888 726 2896 730
rect 2898 732 2906 735
rect 2898 728 2900 732
rect 2904 728 2906 732
rect 2898 726 2906 728
rect 2833 722 2839 723
rect 2833 718 2834 722
rect 2838 718 2839 722
rect 2833 717 2839 718
rect 2901 723 2906 726
rect 2908 723 2913 735
rect 2915 723 2923 735
rect 2933 734 2940 735
rect 2933 730 2934 734
rect 2938 730 2940 734
rect 2933 729 2940 730
rect 2942 732 2950 735
rect 2942 729 2952 732
rect 2944 723 2952 729
rect 2954 723 2959 732
rect 2961 731 2968 732
rect 2961 727 2963 731
rect 2967 727 2968 731
rect 2961 726 2968 727
rect 2961 723 2966 726
rect 2917 722 2923 723
rect 2917 718 2918 722
rect 2922 718 2923 722
rect 2917 717 2923 718
rect 2944 722 2950 723
rect 2944 718 2945 722
rect 2949 718 2950 722
rect 2944 717 2950 718
rect 2584 715 2590 716
rect 2059 709 2066 710
rect 2059 705 2061 709
rect 2065 705 2066 709
rect 2059 704 2066 705
rect 2078 706 2085 707
rect 2039 697 2044 704
rect 1746 690 1755 692
rect 2078 702 2079 706
rect 2083 702 2085 706
rect 2078 701 2085 702
rect 2087 706 2095 707
rect 2087 702 2089 706
rect 2093 702 2095 706
rect 2087 701 2095 702
rect 2097 706 2105 707
rect 2097 702 2099 706
rect 2103 702 2105 706
rect 2097 701 2105 702
rect 2107 706 2114 707
rect 2107 702 2109 706
rect 2113 702 2114 706
rect 2107 701 2114 702
rect 1746 683 1755 688
rect 1746 679 1755 681
rect 1149 666 1160 669
rect 1162 666 1179 669
rect 1189 668 1199 669
rect 1189 664 1191 668
rect 1195 664 1199 668
rect 1189 663 1199 664
rect 1201 663 1220 669
rect 1222 668 1230 669
rect 1222 664 1225 668
rect 1229 664 1230 668
rect 1222 663 1230 664
rect 1243 668 1253 669
rect 1243 664 1245 668
rect 1249 664 1253 668
rect 1243 663 1253 664
rect 1255 663 1274 669
rect 1276 668 1284 669
rect 1276 664 1279 668
rect 1283 664 1284 668
rect 1276 663 1284 664
rect 1299 668 1309 669
rect 1299 664 1301 668
rect 1305 664 1309 668
rect 1299 663 1309 664
rect 1311 663 1330 669
rect 1332 668 1340 669
rect 1332 664 1335 668
rect 1339 664 1340 668
rect 1332 663 1340 664
rect 1353 668 1363 669
rect 1353 664 1355 668
rect 1359 664 1363 668
rect 1353 663 1363 664
rect 1365 663 1384 669
rect 1386 668 1394 669
rect 1627 668 1633 669
rect 1386 664 1389 668
rect 1393 664 1394 668
rect 1386 663 1394 664
rect 1627 664 1628 668
rect 1632 664 1633 668
rect 1627 662 1633 664
rect 1743 678 1761 679
rect 1743 674 1756 678
rect 1760 674 1761 678
rect 1743 673 1761 674
rect 1743 671 1749 673
rect 1627 658 1633 660
rect 1615 657 1633 658
rect 1615 653 1616 657
rect 1620 653 1633 657
rect 1615 652 1633 653
rect 1743 667 1749 669
rect 1743 663 1744 667
rect 1748 663 1749 667
rect 1743 662 1749 663
rect 2794 700 2801 701
rect 2434 698 2441 699
rect 2434 694 2435 698
rect 2439 694 2441 698
rect 2434 693 2441 694
rect 2443 698 2451 699
rect 2443 694 2445 698
rect 2449 694 2451 698
rect 2443 693 2451 694
rect 2453 698 2461 699
rect 2453 694 2455 698
rect 2459 694 2461 698
rect 2453 693 2461 694
rect 2463 698 2470 699
rect 2463 694 2465 698
rect 2469 694 2470 698
rect 2794 696 2795 700
rect 2799 696 2801 700
rect 2794 695 2801 696
rect 2803 700 2811 701
rect 2803 696 2805 700
rect 2809 696 2811 700
rect 2803 695 2811 696
rect 2813 700 2821 701
rect 2813 696 2815 700
rect 2819 696 2821 700
rect 2813 695 2821 696
rect 2823 700 2830 701
rect 2823 696 2825 700
rect 2829 696 2830 700
rect 2823 695 2830 696
rect 2463 693 2470 694
rect 1621 650 1630 652
rect 1621 643 1630 648
rect 1621 639 1630 641
rect 1621 636 1625 639
rect 1624 635 1625 636
rect 1629 635 1630 639
rect 1624 634 1630 635
rect 1743 651 1761 652
rect 1743 647 1756 651
rect 1760 647 1761 651
rect 1743 646 1761 647
rect 1743 644 1755 646
rect 1743 637 1755 642
rect 1743 633 1755 635
rect 1743 629 1746 633
rect 1750 630 1755 633
rect 1750 629 1752 630
rect 1743 627 1752 629
rect 1743 623 1752 625
rect 1743 619 1744 623
rect 1748 619 1752 623
rect 1743 617 1752 619
rect 374 609 379 612
rect 372 608 379 609
rect 372 604 373 608
rect 377 604 379 608
rect 372 603 379 604
rect 381 603 392 612
rect 383 601 392 603
rect 394 601 399 612
rect 401 607 406 612
rect 467 609 472 612
rect 465 608 472 609
rect 401 606 408 607
rect 401 602 403 606
rect 407 602 408 606
rect 465 604 466 608
rect 470 604 472 608
rect 465 603 472 604
rect 474 603 485 612
rect 401 601 408 602
rect 383 596 390 601
rect 476 601 485 603
rect 487 601 492 612
rect 494 607 499 612
rect 554 609 559 612
rect 552 608 559 609
rect 494 606 501 607
rect 494 602 496 606
rect 500 602 501 606
rect 552 604 553 608
rect 557 604 559 608
rect 552 603 559 604
rect 561 603 572 612
rect 494 601 501 602
rect 383 592 384 596
rect 388 592 390 596
rect 383 591 390 592
rect 476 596 483 601
rect 563 601 572 603
rect 574 601 579 612
rect 581 607 586 612
rect 1743 611 1752 615
rect 581 606 588 607
rect 581 602 583 606
rect 587 602 588 606
rect 581 601 588 602
rect 476 592 477 596
rect 481 592 483 596
rect 476 591 483 592
rect 563 596 570 601
rect 1743 607 1747 611
rect 1751 607 1752 611
rect 1743 606 1752 607
rect 1738 601 1747 606
rect 563 592 564 596
rect 568 592 570 596
rect 1738 597 1747 599
rect 1738 593 1739 597
rect 1743 594 1747 597
rect 1743 593 1744 594
rect 1738 592 1744 593
rect 563 591 570 592
rect 1632 590 1638 591
rect 1632 589 1633 590
rect 1629 586 1633 589
rect 1637 586 1638 590
rect 1629 584 1638 586
rect 1593 575 1599 576
rect 1593 571 1594 575
rect 1598 571 1599 575
rect 1593 569 1599 571
rect 1593 565 1599 567
rect 1593 561 1594 565
rect 1598 561 1599 565
rect 1593 559 1599 561
rect 1593 555 1599 557
rect 1593 551 1594 555
rect 1598 551 1599 555
rect 1593 549 1599 551
rect 1593 545 1599 547
rect 1593 541 1594 545
rect 1598 541 1599 545
rect 1629 577 1638 582
rect 1624 576 1633 577
rect 1624 572 1625 576
rect 1629 572 1633 576
rect 1624 568 1633 572
rect 1624 564 1633 566
rect 1624 560 1628 564
rect 1632 560 1633 564
rect 1624 558 1633 560
rect 1743 567 1761 568
rect 1743 563 1756 567
rect 1760 563 1761 567
rect 1743 562 1761 563
rect 1743 560 1755 562
rect 1624 554 1633 556
rect 1624 553 1626 554
rect 1621 550 1626 553
rect 1630 550 1633 554
rect 1621 548 1633 550
rect 1777 558 1783 559
rect 1743 553 1755 558
rect 1621 541 1633 546
rect 1593 540 1599 541
rect 1743 549 1755 551
rect 1743 545 1746 549
rect 1750 546 1755 549
rect 1750 545 1752 546
rect 1743 543 1752 545
rect 1621 537 1633 539
rect 1615 536 1633 537
rect 1615 532 1616 536
rect 1620 532 1633 536
rect 1615 531 1633 532
rect 1743 539 1752 541
rect 1743 535 1744 539
rect 1748 535 1752 539
rect 1743 533 1752 535
rect 186 523 193 524
rect 186 519 188 523
rect 192 519 193 523
rect 186 514 193 519
rect 273 523 280 524
rect 273 519 275 523
rect 279 519 280 523
rect 168 513 175 514
rect 168 509 169 513
rect 173 509 175 513
rect 168 508 175 509
rect 170 503 175 508
rect 177 503 182 514
rect 184 512 193 514
rect 273 514 280 519
rect 366 523 373 524
rect 366 519 368 523
rect 372 519 373 523
rect 255 513 262 514
rect 184 503 195 512
rect 197 511 204 512
rect 197 507 199 511
rect 203 507 204 511
rect 255 509 256 513
rect 260 509 262 513
rect 255 508 262 509
rect 197 506 204 507
rect 197 503 202 506
rect 257 503 262 508
rect 264 503 269 514
rect 271 512 280 514
rect 366 514 373 519
rect 599 525 606 526
rect 599 521 600 525
rect 604 521 606 525
rect 348 513 355 514
rect 271 503 282 512
rect 284 511 291 512
rect 284 507 286 511
rect 290 507 291 511
rect 348 509 349 513
rect 353 509 355 513
rect 348 508 355 509
rect 284 506 291 507
rect 284 503 289 506
rect 350 503 355 508
rect 357 503 362 514
rect 364 512 373 514
rect 599 516 606 521
rect 692 525 699 526
rect 692 521 693 525
rect 697 521 699 525
rect 599 514 608 516
rect 588 513 595 514
rect 364 503 375 512
rect 377 511 384 512
rect 377 507 379 511
rect 383 507 384 511
rect 588 509 589 513
rect 593 509 595 513
rect 588 508 595 509
rect 377 506 384 507
rect 377 503 382 506
rect 590 505 595 508
rect 597 505 608 514
rect 610 505 615 516
rect 617 515 624 516
rect 617 511 619 515
rect 623 511 624 515
rect 692 516 699 521
rect 779 525 786 526
rect 779 521 780 525
rect 784 521 786 525
rect 1743 527 1752 531
rect 692 514 701 516
rect 617 510 624 511
rect 681 513 688 514
rect 617 505 622 510
rect 681 509 682 513
rect 686 509 688 513
rect 681 508 688 509
rect 683 505 688 508
rect 690 505 701 514
rect 703 505 708 516
rect 710 515 717 516
rect 710 511 712 515
rect 716 511 717 515
rect 779 516 786 521
rect 1743 523 1747 527
rect 1751 523 1752 527
rect 1743 522 1752 523
rect 1738 517 1747 522
rect 1777 554 1778 558
rect 1782 554 1783 558
rect 1777 552 1783 554
rect 1777 548 1783 550
rect 1777 544 1778 548
rect 1782 544 1783 548
rect 1777 542 1783 544
rect 1777 538 1783 540
rect 1777 534 1778 538
rect 1782 534 1783 538
rect 1777 532 1783 534
rect 1777 528 1783 530
rect 1777 524 1778 528
rect 1782 524 1783 528
rect 1777 523 1783 524
rect 779 514 788 516
rect 710 510 717 511
rect 768 513 775 514
rect 710 505 715 510
rect 768 509 769 513
rect 773 509 775 513
rect 768 508 775 509
rect 770 505 775 508
rect 777 505 788 514
rect 790 505 795 516
rect 797 515 804 516
rect 797 511 799 515
rect 803 511 804 515
rect 797 510 804 511
rect 797 505 802 510
rect 1738 513 1747 515
rect 1738 509 1739 513
rect 1743 510 1747 513
rect 1743 509 1744 510
rect 1738 508 1744 509
rect 1632 506 1638 507
rect 1632 505 1633 506
rect 1629 502 1633 505
rect 1637 502 1638 506
rect 1629 500 1638 502
rect 1095 465 1106 468
rect 1108 465 1125 468
rect 1629 493 1638 498
rect 1624 492 1633 493
rect 1624 488 1625 492
rect 1629 488 1633 492
rect 1624 484 1633 488
rect 1624 480 1633 482
rect 1624 476 1628 480
rect 1632 476 1633 480
rect 1624 474 1633 476
rect 1624 470 1633 472
rect 1207 469 1217 470
rect 1167 464 1178 467
rect 1180 464 1197 467
rect 1207 465 1209 469
rect 1213 465 1217 469
rect 1207 464 1217 465
rect 1219 464 1238 470
rect 1240 469 1248 470
rect 1240 465 1243 469
rect 1247 465 1248 469
rect 1240 464 1248 465
rect 1261 469 1271 470
rect 1261 465 1263 469
rect 1267 465 1271 469
rect 1261 464 1271 465
rect 1273 464 1292 470
rect 1294 469 1302 470
rect 1294 465 1297 469
rect 1301 465 1302 469
rect 1294 464 1302 465
rect 1317 469 1327 470
rect 1317 465 1319 469
rect 1323 465 1327 469
rect 1317 464 1327 465
rect 1329 464 1348 470
rect 1350 469 1358 470
rect 1350 465 1353 469
rect 1357 465 1358 469
rect 1350 464 1358 465
rect 1371 469 1381 470
rect 1371 465 1373 469
rect 1377 465 1381 469
rect 1371 464 1381 465
rect 1383 464 1402 470
rect 1404 469 1412 470
rect 1624 469 1626 470
rect 1404 465 1407 469
rect 1411 465 1412 469
rect 1404 464 1412 465
rect 1621 466 1626 469
rect 1630 466 1633 470
rect 1621 464 1633 466
rect 1621 457 1633 462
rect 1621 453 1633 455
rect 1615 452 1633 453
rect 90 396 97 397
rect 90 392 91 396
rect 95 392 97 396
rect 90 391 97 392
rect 99 394 107 397
rect 168 401 175 402
rect 168 397 169 401
rect 173 397 175 401
rect 168 396 175 397
rect 99 391 109 394
rect 101 385 109 391
rect 111 385 116 394
rect 118 393 125 394
rect 170 393 175 396
rect 177 397 182 402
rect 252 401 259 402
rect 252 397 253 401
rect 257 397 259 401
rect 177 393 191 397
rect 118 389 120 393
rect 124 389 125 393
rect 118 388 125 389
rect 182 389 183 393
rect 187 389 191 393
rect 182 388 191 389
rect 193 396 201 397
rect 193 392 195 396
rect 199 392 201 396
rect 193 388 201 392
rect 203 394 211 397
rect 203 390 205 394
rect 209 390 211 394
rect 203 388 211 390
rect 118 385 123 388
rect 101 384 107 385
rect 101 380 102 384
rect 106 380 107 384
rect 101 379 107 380
rect 206 385 211 388
rect 213 385 218 397
rect 220 385 228 397
rect 252 396 259 397
rect 254 393 259 396
rect 261 397 266 402
rect 261 393 275 397
rect 266 389 267 393
rect 271 389 275 393
rect 266 388 275 389
rect 277 396 285 397
rect 277 392 279 396
rect 283 392 285 396
rect 277 388 285 392
rect 287 394 295 397
rect 287 390 289 394
rect 293 390 295 394
rect 287 388 295 390
rect 222 384 228 385
rect 222 380 223 384
rect 227 380 228 384
rect 222 379 228 380
rect 290 385 295 388
rect 297 385 302 397
rect 304 385 312 397
rect 322 396 329 397
rect 322 392 323 396
rect 327 392 329 396
rect 322 391 329 392
rect 331 394 339 397
rect 419 398 426 399
rect 419 394 420 398
rect 424 394 426 398
rect 331 391 341 394
rect 333 385 341 391
rect 343 385 348 394
rect 350 393 357 394
rect 419 393 426 394
rect 428 396 436 399
rect 497 403 504 404
rect 497 399 498 403
rect 502 399 504 403
rect 497 398 504 399
rect 428 393 438 396
rect 350 389 352 393
rect 356 389 357 393
rect 350 388 357 389
rect 350 385 355 388
rect 430 387 438 393
rect 440 387 445 396
rect 447 395 454 396
rect 499 395 504 398
rect 506 399 511 404
rect 581 403 588 404
rect 581 399 582 403
rect 586 399 588 403
rect 506 395 520 399
rect 447 391 449 395
rect 453 391 454 395
rect 447 390 454 391
rect 511 391 512 395
rect 516 391 520 395
rect 511 390 520 391
rect 522 398 530 399
rect 522 394 524 398
rect 528 394 530 398
rect 522 390 530 394
rect 532 396 540 399
rect 532 392 534 396
rect 538 392 540 396
rect 532 390 540 392
rect 447 387 452 390
rect 306 384 312 385
rect 306 380 307 384
rect 311 380 312 384
rect 306 379 312 380
rect 333 384 339 385
rect 333 380 334 384
rect 338 380 339 384
rect 430 386 436 387
rect 430 382 431 386
rect 435 382 436 386
rect 430 381 436 382
rect 535 387 540 390
rect 542 387 547 399
rect 549 387 557 399
rect 581 398 588 399
rect 583 395 588 398
rect 590 399 595 404
rect 590 395 604 399
rect 595 391 596 395
rect 600 391 604 395
rect 595 390 604 391
rect 606 398 614 399
rect 606 394 608 398
rect 612 394 614 398
rect 606 390 614 394
rect 616 396 624 399
rect 616 392 618 396
rect 622 392 624 396
rect 616 390 624 392
rect 551 386 557 387
rect 551 382 552 386
rect 556 382 557 386
rect 551 381 557 382
rect 619 387 624 390
rect 626 387 631 399
rect 633 387 641 399
rect 651 398 658 399
rect 651 394 652 398
rect 656 394 658 398
rect 651 393 658 394
rect 660 396 668 399
rect 746 401 753 402
rect 746 397 747 401
rect 751 397 753 401
rect 746 396 753 397
rect 755 399 763 402
rect 1615 448 1616 452
rect 1620 448 1633 452
rect 1615 447 1633 448
rect 1746 464 1752 465
rect 1746 460 1747 464
rect 1751 463 1752 464
rect 1751 460 1755 463
rect 1746 458 1755 460
rect 1746 451 1755 456
rect 2051 452 2058 453
rect 1746 447 1755 449
rect 2051 448 2053 452
rect 2057 448 2058 452
rect 1171 442 1182 445
rect 1184 442 1201 445
rect 1211 444 1221 445
rect 1211 440 1213 444
rect 1217 440 1221 444
rect 1211 439 1221 440
rect 1223 439 1242 445
rect 1244 444 1252 445
rect 1244 440 1247 444
rect 1251 440 1252 444
rect 1244 439 1252 440
rect 1265 444 1275 445
rect 1265 440 1267 444
rect 1271 440 1275 444
rect 1265 439 1275 440
rect 1277 439 1296 445
rect 1298 444 1306 445
rect 1298 440 1301 444
rect 1305 440 1306 444
rect 1298 439 1306 440
rect 1321 444 1331 445
rect 1321 440 1323 444
rect 1327 440 1331 444
rect 1321 439 1331 440
rect 1333 439 1352 445
rect 1354 444 1362 445
rect 1354 440 1357 444
rect 1361 440 1362 444
rect 1354 439 1362 440
rect 1375 444 1385 445
rect 1375 440 1377 444
rect 1381 440 1385 444
rect 1375 439 1385 440
rect 1387 439 1406 445
rect 1408 444 1416 445
rect 1408 440 1411 444
rect 1415 440 1416 444
rect 1408 439 1416 440
rect 1627 436 1633 437
rect 1627 432 1628 436
rect 1632 432 1633 436
rect 1627 430 1633 432
rect 1743 446 1761 447
rect 1743 442 1756 446
rect 1760 442 1761 446
rect 2051 443 2058 448
rect 2138 452 2145 453
rect 2138 448 2140 452
rect 2144 448 2145 452
rect 1743 441 1761 442
rect 2033 442 2040 443
rect 1743 439 1749 441
rect 2033 438 2034 442
rect 2038 438 2040 442
rect 2033 437 2040 438
rect 1627 426 1633 428
rect 1615 425 1633 426
rect 1615 421 1616 425
rect 1620 421 1633 425
rect 1615 420 1633 421
rect 1743 435 1749 437
rect 1743 431 1744 435
rect 1748 431 1749 435
rect 2035 432 2040 437
rect 2042 432 2047 443
rect 2049 441 2058 443
rect 2138 443 2145 448
rect 2231 452 2238 453
rect 2231 448 2233 452
rect 2237 448 2238 452
rect 2120 442 2127 443
rect 2049 432 2060 441
rect 2062 440 2069 441
rect 2062 436 2064 440
rect 2068 436 2069 440
rect 2120 438 2121 442
rect 2125 438 2127 442
rect 2120 437 2127 438
rect 2062 435 2069 436
rect 2062 432 2067 435
rect 2122 432 2127 437
rect 2129 432 2134 443
rect 2136 441 2145 443
rect 2231 443 2238 448
rect 2464 454 2471 455
rect 2464 450 2465 454
rect 2469 450 2471 454
rect 2213 442 2220 443
rect 2136 432 2147 441
rect 2149 440 2156 441
rect 2149 436 2151 440
rect 2155 436 2156 440
rect 2213 438 2214 442
rect 2218 438 2220 442
rect 2213 437 2220 438
rect 2149 435 2156 436
rect 2149 432 2154 435
rect 2215 432 2220 437
rect 2222 432 2227 443
rect 2229 441 2238 443
rect 2464 445 2471 450
rect 2557 454 2564 455
rect 2557 450 2558 454
rect 2562 450 2564 454
rect 2464 443 2473 445
rect 2453 442 2460 443
rect 2229 432 2240 441
rect 2242 440 2249 441
rect 2242 436 2244 440
rect 2248 436 2249 440
rect 2453 438 2454 442
rect 2458 438 2460 442
rect 2453 437 2460 438
rect 2242 435 2249 436
rect 2242 432 2247 435
rect 2455 434 2460 437
rect 2462 434 2473 443
rect 2475 434 2480 445
rect 2482 444 2489 445
rect 2482 440 2484 444
rect 2488 440 2489 444
rect 2557 445 2564 450
rect 2644 454 2651 455
rect 2644 450 2645 454
rect 2649 450 2651 454
rect 2557 443 2566 445
rect 2482 439 2489 440
rect 2546 442 2553 443
rect 2482 434 2487 439
rect 2546 438 2547 442
rect 2551 438 2553 442
rect 2546 437 2553 438
rect 2548 434 2553 437
rect 2555 434 2566 443
rect 2568 434 2573 445
rect 2575 444 2582 445
rect 2575 440 2577 444
rect 2581 440 2582 444
rect 2644 445 2651 450
rect 2644 443 2653 445
rect 2575 439 2582 440
rect 2633 442 2640 443
rect 2575 434 2580 439
rect 2633 438 2634 442
rect 2638 438 2640 442
rect 2633 437 2640 438
rect 2635 434 2640 437
rect 2642 434 2653 443
rect 2655 434 2660 445
rect 2662 444 2669 445
rect 2662 440 2664 444
rect 2668 440 2669 444
rect 2662 439 2669 440
rect 2662 434 2667 439
rect 1743 430 1749 431
rect 824 406 831 407
rect 824 402 825 406
rect 829 402 831 406
rect 824 401 831 402
rect 755 396 765 399
rect 660 393 670 396
rect 662 387 670 393
rect 672 387 677 396
rect 679 395 686 396
rect 679 391 681 395
rect 685 391 686 395
rect 679 390 686 391
rect 757 390 765 396
rect 767 390 772 399
rect 774 398 781 399
rect 826 398 831 401
rect 833 402 838 407
rect 908 406 915 407
rect 908 402 909 406
rect 913 402 915 406
rect 833 398 847 402
rect 774 394 776 398
rect 780 394 781 398
rect 774 393 781 394
rect 838 394 839 398
rect 843 394 847 398
rect 838 393 847 394
rect 849 401 857 402
rect 849 397 851 401
rect 855 397 857 401
rect 849 393 857 397
rect 859 399 867 402
rect 859 395 861 399
rect 865 395 867 399
rect 859 393 867 395
rect 774 390 779 393
rect 679 387 684 390
rect 635 386 641 387
rect 635 382 636 386
rect 640 382 641 386
rect 635 381 641 382
rect 662 386 668 387
rect 662 382 663 386
rect 667 382 668 386
rect 757 389 763 390
rect 757 385 758 389
rect 762 385 763 389
rect 757 384 763 385
rect 862 390 867 393
rect 869 390 874 402
rect 876 390 884 402
rect 908 401 915 402
rect 910 398 915 401
rect 917 402 922 407
rect 917 398 931 402
rect 922 394 923 398
rect 927 394 931 398
rect 922 393 931 394
rect 933 401 941 402
rect 933 397 935 401
rect 939 397 941 401
rect 933 393 941 397
rect 943 399 951 402
rect 943 395 945 399
rect 949 395 951 399
rect 943 393 951 395
rect 878 389 884 390
rect 878 385 879 389
rect 883 385 884 389
rect 878 384 884 385
rect 946 390 951 393
rect 953 390 958 402
rect 960 390 968 402
rect 978 401 985 402
rect 978 397 979 401
rect 983 397 985 401
rect 978 396 985 397
rect 987 399 995 402
rect 1621 418 1630 420
rect 1621 411 1630 416
rect 1621 407 1630 409
rect 1621 404 1625 407
rect 1624 403 1625 404
rect 1629 403 1630 407
rect 1624 402 1630 403
rect 987 396 997 399
rect 989 390 997 396
rect 999 390 1004 399
rect 1006 398 1013 399
rect 1006 394 1008 398
rect 1012 394 1013 398
rect 1006 393 1013 394
rect 1006 390 1011 393
rect 962 389 968 390
rect 962 385 963 389
rect 967 385 968 389
rect 962 384 968 385
rect 989 389 995 390
rect 989 385 990 389
rect 994 385 995 389
rect 989 384 995 385
rect 662 381 668 382
rect 333 379 339 380
rect 839 367 846 368
rect 512 364 519 365
rect 183 362 190 363
rect 183 358 184 362
rect 188 358 190 362
rect 183 357 190 358
rect 192 362 200 363
rect 192 358 194 362
rect 198 358 200 362
rect 192 357 200 358
rect 202 362 210 363
rect 202 358 204 362
rect 208 358 210 362
rect 202 357 210 358
rect 212 362 219 363
rect 212 358 214 362
rect 218 358 219 362
rect 512 360 513 364
rect 517 360 519 364
rect 512 359 519 360
rect 521 364 529 365
rect 521 360 523 364
rect 527 360 529 364
rect 521 359 529 360
rect 531 364 539 365
rect 531 360 533 364
rect 537 360 539 364
rect 531 359 539 360
rect 541 364 548 365
rect 541 360 543 364
rect 547 360 548 364
rect 839 363 840 367
rect 844 363 846 367
rect 839 362 846 363
rect 848 367 856 368
rect 848 363 850 367
rect 854 363 856 367
rect 848 362 856 363
rect 858 367 866 368
rect 858 363 860 367
rect 864 363 866 367
rect 858 362 866 363
rect 868 367 875 368
rect 868 363 870 367
rect 874 363 875 367
rect 868 362 875 363
rect 541 359 548 360
rect 212 357 219 358
rect 1093 320 1104 323
rect 1106 320 1123 323
rect 1462 339 1470 340
rect 1462 336 1463 339
rect 1453 332 1458 336
rect 1451 331 1458 332
rect 1451 327 1452 331
rect 1456 327 1458 331
rect 1451 326 1458 327
rect 1460 335 1463 336
rect 1467 335 1470 339
rect 1460 326 1470 335
rect 1472 338 1479 340
rect 1472 334 1474 338
rect 1478 334 1479 338
rect 1472 331 1479 334
rect 1472 327 1474 331
rect 1478 327 1479 331
rect 1472 326 1479 327
rect 1738 340 1744 341
rect 1738 336 1739 340
rect 1743 339 1744 340
rect 1743 336 1747 339
rect 1738 334 1747 336
rect 1205 324 1215 325
rect 1165 319 1176 322
rect 1178 319 1195 322
rect 1205 320 1207 324
rect 1211 320 1215 324
rect 1205 319 1215 320
rect 1217 319 1236 325
rect 1238 324 1246 325
rect 1238 320 1241 324
rect 1245 320 1246 324
rect 1238 319 1246 320
rect 1259 324 1269 325
rect 1259 320 1261 324
rect 1265 320 1269 324
rect 1259 319 1269 320
rect 1271 319 1290 325
rect 1292 324 1300 325
rect 1292 320 1295 324
rect 1299 320 1300 324
rect 1292 319 1300 320
rect 1315 324 1325 325
rect 1315 320 1317 324
rect 1321 320 1325 324
rect 1315 319 1325 320
rect 1327 319 1346 325
rect 1348 324 1356 325
rect 1348 320 1351 324
rect 1355 320 1356 324
rect 1348 319 1356 320
rect 1369 324 1379 325
rect 1369 320 1371 324
rect 1375 320 1379 324
rect 1369 319 1379 320
rect 1381 319 1400 325
rect 1402 324 1410 325
rect 1402 320 1405 324
rect 1409 320 1410 324
rect 1402 319 1410 320
rect 1738 327 1747 332
rect 1955 325 1962 326
rect 1738 323 1747 325
rect 89 250 96 251
rect 89 246 90 250
rect 94 246 96 250
rect 89 245 96 246
rect 98 248 106 251
rect 167 255 174 256
rect 167 251 168 255
rect 172 251 174 255
rect 167 250 174 251
rect 98 245 108 248
rect 100 239 108 245
rect 110 239 115 248
rect 117 247 124 248
rect 169 247 174 250
rect 176 251 181 256
rect 251 255 258 256
rect 251 251 252 255
rect 256 251 258 255
rect 176 247 190 251
rect 117 243 119 247
rect 123 243 124 247
rect 117 242 124 243
rect 181 243 182 247
rect 186 243 190 247
rect 181 242 190 243
rect 192 250 200 251
rect 192 246 194 250
rect 198 246 200 250
rect 192 242 200 246
rect 202 248 210 251
rect 202 244 204 248
rect 208 244 210 248
rect 202 242 210 244
rect 117 239 122 242
rect 100 238 106 239
rect 100 234 101 238
rect 105 234 106 238
rect 100 233 106 234
rect 205 239 210 242
rect 212 239 217 251
rect 219 239 227 251
rect 251 250 258 251
rect 253 247 258 250
rect 260 251 265 256
rect 260 247 274 251
rect 265 243 266 247
rect 270 243 274 247
rect 265 242 274 243
rect 276 250 284 251
rect 276 246 278 250
rect 282 246 284 250
rect 276 242 284 246
rect 286 248 294 251
rect 286 244 288 248
rect 292 244 294 248
rect 286 242 294 244
rect 221 238 227 239
rect 221 234 222 238
rect 226 234 227 238
rect 221 233 227 234
rect 289 239 294 242
rect 296 239 301 251
rect 303 239 311 251
rect 321 250 328 251
rect 321 246 322 250
rect 326 246 328 250
rect 321 245 328 246
rect 330 248 338 251
rect 418 252 425 253
rect 418 248 419 252
rect 423 248 425 252
rect 330 245 340 248
rect 332 239 340 245
rect 342 239 347 248
rect 349 247 356 248
rect 418 247 425 248
rect 427 250 435 253
rect 496 257 503 258
rect 496 253 497 257
rect 501 253 503 257
rect 496 252 503 253
rect 427 247 437 250
rect 349 243 351 247
rect 355 243 356 247
rect 349 242 356 243
rect 349 239 354 242
rect 429 241 437 247
rect 439 241 444 250
rect 446 249 453 250
rect 498 249 503 252
rect 505 253 510 258
rect 580 257 587 258
rect 580 253 581 257
rect 585 253 587 257
rect 505 249 519 253
rect 446 245 448 249
rect 452 245 453 249
rect 446 244 453 245
rect 510 245 511 249
rect 515 245 519 249
rect 510 244 519 245
rect 521 252 529 253
rect 521 248 523 252
rect 527 248 529 252
rect 521 244 529 248
rect 531 250 539 253
rect 531 246 533 250
rect 537 246 539 250
rect 531 244 539 246
rect 446 241 451 244
rect 305 238 311 239
rect 305 234 306 238
rect 310 234 311 238
rect 305 233 311 234
rect 332 238 338 239
rect 332 234 333 238
rect 337 234 338 238
rect 429 240 435 241
rect 429 236 430 240
rect 434 236 435 240
rect 429 235 435 236
rect 534 241 539 244
rect 541 241 546 253
rect 548 241 556 253
rect 580 252 587 253
rect 582 249 587 252
rect 589 253 594 258
rect 589 249 603 253
rect 594 245 595 249
rect 599 245 603 249
rect 594 244 603 245
rect 605 252 613 253
rect 605 248 607 252
rect 611 248 613 252
rect 605 244 613 248
rect 615 250 623 253
rect 615 246 617 250
rect 621 246 623 250
rect 615 244 623 246
rect 550 240 556 241
rect 550 236 551 240
rect 555 236 556 240
rect 550 235 556 236
rect 618 241 623 244
rect 625 241 630 253
rect 632 241 640 253
rect 650 252 657 253
rect 650 248 651 252
rect 655 248 657 252
rect 650 247 657 248
rect 659 250 667 253
rect 745 255 752 256
rect 745 251 746 255
rect 750 251 752 255
rect 745 250 752 251
rect 754 253 762 256
rect 1169 297 1180 300
rect 1182 297 1199 300
rect 1209 299 1219 300
rect 1209 295 1211 299
rect 1215 295 1219 299
rect 1209 294 1219 295
rect 1221 294 1240 300
rect 1242 299 1250 300
rect 1242 295 1245 299
rect 1249 295 1250 299
rect 1242 294 1250 295
rect 1263 299 1273 300
rect 1263 295 1265 299
rect 1269 295 1273 299
rect 1263 294 1273 295
rect 1275 294 1294 300
rect 1296 299 1304 300
rect 1296 295 1299 299
rect 1303 295 1304 299
rect 1296 294 1304 295
rect 1319 299 1329 300
rect 1319 295 1321 299
rect 1325 295 1329 299
rect 1319 294 1329 295
rect 1331 294 1350 300
rect 1352 299 1360 300
rect 1352 295 1355 299
rect 1359 295 1360 299
rect 1352 294 1360 295
rect 1373 299 1383 300
rect 1373 295 1375 299
rect 1379 295 1383 299
rect 1373 294 1383 295
rect 1385 294 1404 300
rect 1406 299 1414 300
rect 1406 295 1409 299
rect 1413 295 1414 299
rect 1406 294 1414 295
rect 1735 322 1753 323
rect 1735 318 1748 322
rect 1752 318 1753 322
rect 1955 321 1956 325
rect 1960 321 1962 325
rect 1955 320 1962 321
rect 1964 323 1972 326
rect 2033 330 2040 331
rect 2033 326 2034 330
rect 2038 326 2040 330
rect 2033 325 2040 326
rect 1964 320 1974 323
rect 1735 317 1753 318
rect 1735 315 1741 317
rect 1966 314 1974 320
rect 1976 314 1981 323
rect 1983 322 1990 323
rect 2035 322 2040 325
rect 2042 326 2047 331
rect 2117 330 2124 331
rect 2117 326 2118 330
rect 2122 326 2124 330
rect 2042 322 2056 326
rect 1983 318 1985 322
rect 1989 318 1990 322
rect 1983 317 1990 318
rect 2047 318 2048 322
rect 2052 318 2056 322
rect 2047 317 2056 318
rect 2058 325 2066 326
rect 2058 321 2060 325
rect 2064 321 2066 325
rect 2058 317 2066 321
rect 2068 323 2076 326
rect 2068 319 2070 323
rect 2074 319 2076 323
rect 2068 317 2076 319
rect 1983 314 1988 317
rect 1735 311 1741 313
rect 1735 307 1736 311
rect 1740 307 1741 311
rect 1966 313 1972 314
rect 1966 309 1967 313
rect 1971 309 1972 313
rect 1966 308 1972 309
rect 2071 314 2076 317
rect 2078 314 2083 326
rect 2085 314 2093 326
rect 2117 325 2124 326
rect 2119 322 2124 325
rect 2126 326 2131 331
rect 2126 322 2140 326
rect 2131 318 2132 322
rect 2136 318 2140 322
rect 2131 317 2140 318
rect 2142 325 2150 326
rect 2142 321 2144 325
rect 2148 321 2150 325
rect 2142 317 2150 321
rect 2152 323 2160 326
rect 2152 319 2154 323
rect 2158 319 2160 323
rect 2152 317 2160 319
rect 2087 313 2093 314
rect 2087 309 2088 313
rect 2092 309 2093 313
rect 2087 308 2093 309
rect 2155 314 2160 317
rect 2162 314 2167 326
rect 2169 314 2177 326
rect 2187 325 2194 326
rect 2187 321 2188 325
rect 2192 321 2194 325
rect 2187 320 2194 321
rect 2196 323 2204 326
rect 2284 327 2291 328
rect 2284 323 2285 327
rect 2289 323 2291 327
rect 2196 320 2206 323
rect 2198 314 2206 320
rect 2208 314 2213 323
rect 2215 322 2222 323
rect 2284 322 2291 323
rect 2293 325 2301 328
rect 2362 332 2369 333
rect 2362 328 2363 332
rect 2367 328 2369 332
rect 2362 327 2369 328
rect 2293 322 2303 325
rect 2215 318 2217 322
rect 2221 318 2222 322
rect 2215 317 2222 318
rect 2215 314 2220 317
rect 2295 316 2303 322
rect 2305 316 2310 325
rect 2312 324 2319 325
rect 2364 324 2369 327
rect 2371 328 2376 333
rect 2446 332 2453 333
rect 2446 328 2447 332
rect 2451 328 2453 332
rect 2371 324 2385 328
rect 2312 320 2314 324
rect 2318 320 2319 324
rect 2312 319 2319 320
rect 2376 320 2377 324
rect 2381 320 2385 324
rect 2376 319 2385 320
rect 2387 327 2395 328
rect 2387 323 2389 327
rect 2393 323 2395 327
rect 2387 319 2395 323
rect 2397 325 2405 328
rect 2397 321 2399 325
rect 2403 321 2405 325
rect 2397 319 2405 321
rect 2312 316 2317 319
rect 2171 313 2177 314
rect 2171 309 2172 313
rect 2176 309 2177 313
rect 2171 308 2177 309
rect 2198 313 2204 314
rect 2198 309 2199 313
rect 2203 309 2204 313
rect 2295 315 2301 316
rect 2295 311 2296 315
rect 2300 311 2301 315
rect 2295 310 2301 311
rect 2400 316 2405 319
rect 2407 316 2412 328
rect 2414 316 2422 328
rect 2446 327 2453 328
rect 2448 324 2453 327
rect 2455 328 2460 333
rect 2455 324 2469 328
rect 2460 320 2461 324
rect 2465 320 2469 324
rect 2460 319 2469 320
rect 2471 327 2479 328
rect 2471 323 2473 327
rect 2477 323 2479 327
rect 2471 319 2479 323
rect 2481 325 2489 328
rect 2481 321 2483 325
rect 2487 321 2489 325
rect 2481 319 2489 321
rect 2416 315 2422 316
rect 2416 311 2417 315
rect 2421 311 2422 315
rect 2416 310 2422 311
rect 2484 316 2489 319
rect 2491 316 2496 328
rect 2498 316 2506 328
rect 2516 327 2523 328
rect 2516 323 2517 327
rect 2521 323 2523 327
rect 2516 322 2523 323
rect 2525 325 2533 328
rect 2611 330 2618 331
rect 2611 326 2612 330
rect 2616 326 2618 330
rect 2611 325 2618 326
rect 2620 328 2628 331
rect 2689 335 2696 336
rect 2689 331 2690 335
rect 2694 331 2696 335
rect 2689 330 2696 331
rect 2620 325 2630 328
rect 2525 322 2535 325
rect 2527 316 2535 322
rect 2537 316 2542 325
rect 2544 324 2551 325
rect 2544 320 2546 324
rect 2550 320 2551 324
rect 2544 319 2551 320
rect 2622 319 2630 325
rect 2632 319 2637 328
rect 2639 327 2646 328
rect 2691 327 2696 330
rect 2698 331 2703 336
rect 2773 335 2780 336
rect 2773 331 2774 335
rect 2778 331 2780 335
rect 2698 327 2712 331
rect 2639 323 2641 327
rect 2645 323 2646 327
rect 2639 322 2646 323
rect 2703 323 2704 327
rect 2708 323 2712 327
rect 2703 322 2712 323
rect 2714 330 2722 331
rect 2714 326 2716 330
rect 2720 326 2722 330
rect 2714 322 2722 326
rect 2724 328 2732 331
rect 2724 324 2726 328
rect 2730 324 2732 328
rect 2724 322 2732 324
rect 2639 319 2644 322
rect 2544 316 2549 319
rect 2500 315 2506 316
rect 2500 311 2501 315
rect 2505 311 2506 315
rect 2500 310 2506 311
rect 2527 315 2533 316
rect 2527 311 2528 315
rect 2532 311 2533 315
rect 2622 318 2628 319
rect 2622 314 2623 318
rect 2627 314 2628 318
rect 2622 313 2628 314
rect 2727 319 2732 322
rect 2734 319 2739 331
rect 2741 319 2749 331
rect 2773 330 2780 331
rect 2775 327 2780 330
rect 2782 331 2787 336
rect 2782 327 2796 331
rect 2787 323 2788 327
rect 2792 323 2796 327
rect 2787 322 2796 323
rect 2798 330 2806 331
rect 2798 326 2800 330
rect 2804 326 2806 330
rect 2798 322 2806 326
rect 2808 328 2816 331
rect 2808 324 2810 328
rect 2814 324 2816 328
rect 2808 322 2816 324
rect 2743 318 2749 319
rect 2743 314 2744 318
rect 2748 314 2749 318
rect 2743 313 2749 314
rect 2811 319 2816 322
rect 2818 319 2823 331
rect 2825 319 2833 331
rect 2843 330 2850 331
rect 2843 326 2844 330
rect 2848 326 2850 330
rect 2843 325 2850 326
rect 2852 328 2860 331
rect 2852 325 2862 328
rect 2854 319 2862 325
rect 2864 319 2869 328
rect 2871 327 2878 328
rect 2871 323 2873 327
rect 2877 323 2878 327
rect 2871 322 2878 323
rect 2871 319 2876 322
rect 2827 318 2833 319
rect 2827 314 2828 318
rect 2832 314 2833 318
rect 2827 313 2833 314
rect 2854 318 2860 319
rect 2854 314 2855 318
rect 2859 314 2860 318
rect 2854 313 2860 314
rect 2527 310 2533 311
rect 2198 308 2204 309
rect 1735 306 1741 307
rect 1735 295 1753 296
rect 1735 291 1748 295
rect 1752 291 1753 295
rect 2704 296 2711 297
rect 2377 293 2384 294
rect 1735 290 1753 291
rect 2048 291 2055 292
rect 1735 288 1747 290
rect 2048 287 2049 291
rect 2053 287 2055 291
rect 2048 286 2055 287
rect 2057 291 2065 292
rect 2057 287 2059 291
rect 2063 287 2065 291
rect 2057 286 2065 287
rect 2067 291 2075 292
rect 2067 287 2069 291
rect 2073 287 2075 291
rect 2067 286 2075 287
rect 2077 291 2084 292
rect 2077 287 2079 291
rect 2083 287 2084 291
rect 2377 289 2378 293
rect 2382 289 2384 293
rect 2377 288 2384 289
rect 2386 293 2394 294
rect 2386 289 2388 293
rect 2392 289 2394 293
rect 2386 288 2394 289
rect 2396 293 2404 294
rect 2396 289 2398 293
rect 2402 289 2404 293
rect 2396 288 2404 289
rect 2406 293 2413 294
rect 2406 289 2408 293
rect 2412 289 2413 293
rect 2704 292 2705 296
rect 2709 292 2711 296
rect 2704 291 2711 292
rect 2713 296 2721 297
rect 2713 292 2715 296
rect 2719 292 2721 296
rect 2713 291 2721 292
rect 2723 296 2731 297
rect 2723 292 2725 296
rect 2729 292 2731 296
rect 2723 291 2731 292
rect 2733 296 2740 297
rect 2733 292 2735 296
rect 2739 292 2740 296
rect 2733 291 2740 292
rect 2406 288 2413 289
rect 2077 286 2084 287
rect 1735 281 1747 286
rect 823 260 830 261
rect 823 256 824 260
rect 828 256 830 260
rect 823 255 830 256
rect 754 250 764 253
rect 659 247 669 250
rect 661 241 669 247
rect 671 241 676 250
rect 678 249 685 250
rect 678 245 680 249
rect 684 245 685 249
rect 678 244 685 245
rect 756 244 764 250
rect 766 244 771 253
rect 773 252 780 253
rect 825 252 830 255
rect 832 256 837 261
rect 907 260 914 261
rect 907 256 908 260
rect 912 256 914 260
rect 832 252 846 256
rect 773 248 775 252
rect 779 248 780 252
rect 773 247 780 248
rect 837 248 838 252
rect 842 248 846 252
rect 837 247 846 248
rect 848 255 856 256
rect 848 251 850 255
rect 854 251 856 255
rect 848 247 856 251
rect 858 253 866 256
rect 858 249 860 253
rect 864 249 866 253
rect 858 247 866 249
rect 773 244 778 247
rect 678 241 683 244
rect 634 240 640 241
rect 634 236 635 240
rect 639 236 640 240
rect 634 235 640 236
rect 661 240 667 241
rect 661 236 662 240
rect 666 236 667 240
rect 756 243 762 244
rect 756 239 757 243
rect 761 239 762 243
rect 756 238 762 239
rect 861 244 866 247
rect 868 244 873 256
rect 875 244 883 256
rect 907 255 914 256
rect 909 252 914 255
rect 916 256 921 261
rect 916 252 930 256
rect 921 248 922 252
rect 926 248 930 252
rect 921 247 930 248
rect 932 255 940 256
rect 932 251 934 255
rect 938 251 940 255
rect 932 247 940 251
rect 942 253 950 256
rect 942 249 944 253
rect 948 249 950 253
rect 942 247 950 249
rect 877 243 883 244
rect 877 239 878 243
rect 882 239 883 243
rect 877 238 883 239
rect 945 244 950 247
rect 952 244 957 256
rect 959 244 967 256
rect 977 255 984 256
rect 977 251 978 255
rect 982 251 984 255
rect 977 250 984 251
rect 986 253 994 256
rect 1735 277 1747 279
rect 1735 273 1738 277
rect 1742 274 1747 277
rect 1742 273 1744 274
rect 1735 271 1744 273
rect 1735 267 1744 269
rect 1735 263 1736 267
rect 1740 263 1744 267
rect 1735 261 1744 263
rect 986 250 996 253
rect 988 244 996 250
rect 998 244 1003 253
rect 1005 252 1012 253
rect 1005 248 1007 252
rect 1011 248 1012 252
rect 1005 247 1012 248
rect 1005 244 1010 247
rect 961 243 967 244
rect 961 239 962 243
rect 966 239 967 243
rect 961 238 967 239
rect 988 243 994 244
rect 988 239 989 243
rect 993 239 994 243
rect 988 238 994 239
rect 661 235 667 236
rect 332 233 338 234
rect 838 221 845 222
rect 511 218 518 219
rect 182 216 189 217
rect 182 212 183 216
rect 187 212 189 216
rect 182 211 189 212
rect 191 216 199 217
rect 191 212 193 216
rect 197 212 199 216
rect 191 211 199 212
rect 201 216 209 217
rect 201 212 203 216
rect 207 212 209 216
rect 201 211 209 212
rect 211 216 218 217
rect 211 212 213 216
rect 217 212 218 216
rect 511 214 512 218
rect 516 214 518 218
rect 511 213 518 214
rect 520 218 528 219
rect 520 214 522 218
rect 526 214 528 218
rect 520 213 528 214
rect 530 218 538 219
rect 530 214 532 218
rect 536 214 538 218
rect 530 213 538 214
rect 540 218 547 219
rect 540 214 542 218
rect 546 214 547 218
rect 838 217 839 221
rect 843 217 845 221
rect 838 216 845 217
rect 847 221 855 222
rect 847 217 849 221
rect 853 217 855 221
rect 847 216 855 217
rect 857 221 865 222
rect 857 217 859 221
rect 863 217 865 221
rect 857 216 865 217
rect 867 221 874 222
rect 867 217 869 221
rect 873 217 874 221
rect 867 216 874 217
rect 540 213 547 214
rect 211 211 218 212
rect 1735 255 1744 259
rect 1735 251 1739 255
rect 1743 251 1744 255
rect 1735 250 1744 251
rect 1730 245 1739 250
rect 1730 241 1739 243
rect 1730 237 1731 241
rect 1735 238 1739 241
rect 1735 237 1736 238
rect 1730 236 1736 237
rect 1453 212 1460 213
rect 1453 208 1454 212
rect 1458 208 1460 212
rect 1453 207 1460 208
rect 1455 203 1460 207
rect 1462 204 1472 213
rect 1462 203 1465 204
rect 1464 200 1465 203
rect 1469 200 1472 204
rect 1464 199 1472 200
rect 1474 212 1481 213
rect 1474 208 1476 212
rect 1480 208 1481 212
rect 1474 205 1481 208
rect 1735 211 1753 212
rect 1735 207 1748 211
rect 1752 207 1753 211
rect 1735 206 1753 207
rect 1474 201 1476 205
rect 1480 201 1481 205
rect 1735 204 1747 206
rect 1474 199 1481 201
rect 1094 178 1105 181
rect 1107 178 1124 181
rect 1769 202 1775 203
rect 1735 197 1747 202
rect 1735 193 1747 195
rect 1735 189 1738 193
rect 1742 190 1747 193
rect 1742 189 1744 190
rect 1735 187 1744 189
rect 1206 182 1216 183
rect 1166 177 1177 180
rect 1179 177 1196 180
rect 1206 178 1208 182
rect 1212 178 1216 182
rect 1206 177 1216 178
rect 1218 177 1237 183
rect 1239 182 1247 183
rect 1239 178 1242 182
rect 1246 178 1247 182
rect 1239 177 1247 178
rect 1260 182 1270 183
rect 1260 178 1262 182
rect 1266 178 1270 182
rect 1260 177 1270 178
rect 1272 177 1291 183
rect 1293 182 1301 183
rect 1293 178 1296 182
rect 1300 178 1301 182
rect 1293 177 1301 178
rect 1316 182 1326 183
rect 1316 178 1318 182
rect 1322 178 1326 182
rect 1316 177 1326 178
rect 1328 177 1347 183
rect 1349 182 1357 183
rect 1349 178 1352 182
rect 1356 178 1357 182
rect 1349 177 1357 178
rect 1370 182 1380 183
rect 1370 178 1372 182
rect 1376 178 1380 182
rect 1370 177 1380 178
rect 1382 177 1401 183
rect 1403 182 1411 183
rect 1403 178 1406 182
rect 1410 178 1411 182
rect 1403 177 1411 178
rect 1735 183 1744 185
rect 1735 179 1736 183
rect 1740 179 1744 183
rect 1735 177 1744 179
rect 1735 171 1744 175
rect 1170 155 1181 158
rect 1183 155 1200 158
rect 1210 157 1220 158
rect 1210 153 1212 157
rect 1216 153 1220 157
rect 1210 152 1220 153
rect 1222 152 1241 158
rect 1243 157 1251 158
rect 1243 153 1246 157
rect 1250 153 1251 157
rect 1243 152 1251 153
rect 1264 157 1274 158
rect 1264 153 1266 157
rect 1270 153 1274 157
rect 1264 152 1274 153
rect 1276 152 1295 158
rect 1297 157 1305 158
rect 1297 153 1300 157
rect 1304 153 1305 157
rect 1297 152 1305 153
rect 1320 157 1330 158
rect 1320 153 1322 157
rect 1326 153 1330 157
rect 1320 152 1330 153
rect 1332 152 1351 158
rect 1353 157 1361 158
rect 1353 153 1356 157
rect 1360 153 1361 157
rect 1353 152 1361 153
rect 1374 157 1384 158
rect 1374 153 1376 157
rect 1380 153 1384 157
rect 1374 152 1384 153
rect 1386 152 1405 158
rect 1407 157 1415 158
rect 1466 160 1474 161
rect 1466 157 1467 160
rect 1407 153 1410 157
rect 1414 153 1415 157
rect 1457 153 1462 157
rect 1407 152 1415 153
rect 1455 152 1462 153
rect 1455 148 1456 152
rect 1460 148 1462 152
rect 1455 147 1462 148
rect 1464 156 1467 157
rect 1471 156 1474 160
rect 1464 147 1474 156
rect 1476 159 1483 161
rect 1735 167 1739 171
rect 1743 167 1744 171
rect 1735 166 1744 167
rect 1730 161 1739 166
rect 1769 198 1770 202
rect 1774 198 1775 202
rect 1769 196 1775 198
rect 1769 192 1775 194
rect 1769 188 1770 192
rect 1774 188 1775 192
rect 1769 186 1775 188
rect 1769 182 1775 184
rect 1769 178 1770 182
rect 1774 178 1775 182
rect 1769 176 1775 178
rect 1954 179 1961 180
rect 1769 172 1775 174
rect 1769 168 1770 172
rect 1774 168 1775 172
rect 1954 175 1955 179
rect 1959 175 1961 179
rect 1954 174 1961 175
rect 1963 177 1971 180
rect 2032 184 2039 185
rect 2032 180 2033 184
rect 2037 180 2039 184
rect 2032 179 2039 180
rect 1963 174 1973 177
rect 1769 167 1775 168
rect 1965 168 1973 174
rect 1975 168 1980 177
rect 1982 176 1989 177
rect 2034 176 2039 179
rect 2041 180 2046 185
rect 2116 184 2123 185
rect 2116 180 2117 184
rect 2121 180 2123 184
rect 2041 176 2055 180
rect 1982 172 1984 176
rect 1988 172 1989 176
rect 1982 171 1989 172
rect 2046 172 2047 176
rect 2051 172 2055 176
rect 2046 171 2055 172
rect 2057 179 2065 180
rect 2057 175 2059 179
rect 2063 175 2065 179
rect 2057 171 2065 175
rect 2067 177 2075 180
rect 2067 173 2069 177
rect 2073 173 2075 177
rect 2067 171 2075 173
rect 1982 168 1987 171
rect 1965 167 1971 168
rect 1965 163 1966 167
rect 1970 163 1971 167
rect 1965 162 1971 163
rect 2070 168 2075 171
rect 2077 168 2082 180
rect 2084 168 2092 180
rect 2116 179 2123 180
rect 2118 176 2123 179
rect 2125 180 2130 185
rect 2125 176 2139 180
rect 2130 172 2131 176
rect 2135 172 2139 176
rect 2130 171 2139 172
rect 2141 179 2149 180
rect 2141 175 2143 179
rect 2147 175 2149 179
rect 2141 171 2149 175
rect 2151 177 2159 180
rect 2151 173 2153 177
rect 2157 173 2159 177
rect 2151 171 2159 173
rect 2086 167 2092 168
rect 2086 163 2087 167
rect 2091 163 2092 167
rect 2086 162 2092 163
rect 2154 168 2159 171
rect 2161 168 2166 180
rect 2168 168 2176 180
rect 2186 179 2193 180
rect 2186 175 2187 179
rect 2191 175 2193 179
rect 2186 174 2193 175
rect 2195 177 2203 180
rect 2283 181 2290 182
rect 2283 177 2284 181
rect 2288 177 2290 181
rect 2195 174 2205 177
rect 2197 168 2205 174
rect 2207 168 2212 177
rect 2214 176 2221 177
rect 2283 176 2290 177
rect 2292 179 2300 182
rect 2361 186 2368 187
rect 2361 182 2362 186
rect 2366 182 2368 186
rect 2361 181 2368 182
rect 2292 176 2302 179
rect 2214 172 2216 176
rect 2220 172 2221 176
rect 2214 171 2221 172
rect 2214 168 2219 171
rect 2294 170 2302 176
rect 2304 170 2309 179
rect 2311 178 2318 179
rect 2363 178 2368 181
rect 2370 182 2375 187
rect 2445 186 2452 187
rect 2445 182 2446 186
rect 2450 182 2452 186
rect 2370 178 2384 182
rect 2311 174 2313 178
rect 2317 174 2318 178
rect 2311 173 2318 174
rect 2375 174 2376 178
rect 2380 174 2384 178
rect 2375 173 2384 174
rect 2386 181 2394 182
rect 2386 177 2388 181
rect 2392 177 2394 181
rect 2386 173 2394 177
rect 2396 179 2404 182
rect 2396 175 2398 179
rect 2402 175 2404 179
rect 2396 173 2404 175
rect 2311 170 2316 173
rect 2170 167 2176 168
rect 2170 163 2171 167
rect 2175 163 2176 167
rect 2170 162 2176 163
rect 2197 167 2203 168
rect 2197 163 2198 167
rect 2202 163 2203 167
rect 2294 169 2300 170
rect 2294 165 2295 169
rect 2299 165 2300 169
rect 2294 164 2300 165
rect 2399 170 2404 173
rect 2406 170 2411 182
rect 2413 170 2421 182
rect 2445 181 2452 182
rect 2447 178 2452 181
rect 2454 182 2459 187
rect 2454 178 2468 182
rect 2459 174 2460 178
rect 2464 174 2468 178
rect 2459 173 2468 174
rect 2470 181 2478 182
rect 2470 177 2472 181
rect 2476 177 2478 181
rect 2470 173 2478 177
rect 2480 179 2488 182
rect 2480 175 2482 179
rect 2486 175 2488 179
rect 2480 173 2488 175
rect 2415 169 2421 170
rect 2415 165 2416 169
rect 2420 165 2421 169
rect 2415 164 2421 165
rect 2483 170 2488 173
rect 2490 170 2495 182
rect 2497 170 2505 182
rect 2515 181 2522 182
rect 2515 177 2516 181
rect 2520 177 2522 181
rect 2515 176 2522 177
rect 2524 179 2532 182
rect 2610 184 2617 185
rect 2610 180 2611 184
rect 2615 180 2617 184
rect 2610 179 2617 180
rect 2619 182 2627 185
rect 2688 189 2695 190
rect 2688 185 2689 189
rect 2693 185 2695 189
rect 2688 184 2695 185
rect 2619 179 2629 182
rect 2524 176 2534 179
rect 2526 170 2534 176
rect 2536 170 2541 179
rect 2543 178 2550 179
rect 2543 174 2545 178
rect 2549 174 2550 178
rect 2543 173 2550 174
rect 2621 173 2629 179
rect 2631 173 2636 182
rect 2638 181 2645 182
rect 2690 181 2695 184
rect 2697 185 2702 190
rect 2772 189 2779 190
rect 2772 185 2773 189
rect 2777 185 2779 189
rect 2697 181 2711 185
rect 2638 177 2640 181
rect 2644 177 2645 181
rect 2638 176 2645 177
rect 2702 177 2703 181
rect 2707 177 2711 181
rect 2702 176 2711 177
rect 2713 184 2721 185
rect 2713 180 2715 184
rect 2719 180 2721 184
rect 2713 176 2721 180
rect 2723 182 2731 185
rect 2723 178 2725 182
rect 2729 178 2731 182
rect 2723 176 2731 178
rect 2638 173 2643 176
rect 2543 170 2548 173
rect 2499 169 2505 170
rect 2499 165 2500 169
rect 2504 165 2505 169
rect 2499 164 2505 165
rect 2526 169 2532 170
rect 2526 165 2527 169
rect 2531 165 2532 169
rect 2621 172 2627 173
rect 2621 168 2622 172
rect 2626 168 2627 172
rect 2621 167 2627 168
rect 2726 173 2731 176
rect 2733 173 2738 185
rect 2740 173 2748 185
rect 2772 184 2779 185
rect 2774 181 2779 184
rect 2781 185 2786 190
rect 2781 181 2795 185
rect 2786 177 2787 181
rect 2791 177 2795 181
rect 2786 176 2795 177
rect 2797 184 2805 185
rect 2797 180 2799 184
rect 2803 180 2805 184
rect 2797 176 2805 180
rect 2807 182 2815 185
rect 2807 178 2809 182
rect 2813 178 2815 182
rect 2807 176 2815 178
rect 2742 172 2748 173
rect 2742 168 2743 172
rect 2747 168 2748 172
rect 2742 167 2748 168
rect 2810 173 2815 176
rect 2817 173 2822 185
rect 2824 173 2832 185
rect 2842 184 2849 185
rect 2842 180 2843 184
rect 2847 180 2849 184
rect 2842 179 2849 180
rect 2851 182 2859 185
rect 2851 179 2861 182
rect 2853 173 2861 179
rect 2863 173 2868 182
rect 2870 181 2877 182
rect 2870 177 2872 181
rect 2876 177 2877 181
rect 2870 176 2877 177
rect 2870 173 2875 176
rect 2826 172 2832 173
rect 2826 168 2827 172
rect 2831 168 2832 172
rect 2826 167 2832 168
rect 2853 172 2859 173
rect 2853 168 2854 172
rect 2858 168 2859 172
rect 2853 167 2859 168
rect 2526 164 2532 165
rect 2197 162 2203 163
rect 1476 155 1478 159
rect 1482 155 1483 159
rect 1476 152 1483 155
rect 1730 157 1739 159
rect 1730 153 1731 157
rect 1735 154 1739 157
rect 1735 153 1736 154
rect 1766 154 1772 155
rect 1766 153 1767 154
rect 1730 152 1736 153
rect 1476 148 1478 152
rect 1482 148 1483 152
rect 1759 150 1767 153
rect 1771 150 1772 154
rect 1759 148 1772 150
rect 1476 147 1483 148
rect 1759 144 1772 146
rect 1759 141 1763 144
rect 1762 140 1763 141
rect 1767 140 1772 144
rect 2703 150 2710 151
rect 2376 147 2383 148
rect 1762 138 1772 140
rect 385 103 390 106
rect 383 102 390 103
rect 383 98 384 102
rect 388 98 390 102
rect 383 97 390 98
rect 392 97 403 106
rect 394 95 403 97
rect 405 95 410 106
rect 412 101 417 106
rect 478 103 483 106
rect 476 102 483 103
rect 412 100 419 101
rect 412 96 414 100
rect 418 96 419 100
rect 476 98 477 102
rect 481 98 483 102
rect 476 97 483 98
rect 485 97 496 106
rect 412 95 419 96
rect 394 90 401 95
rect 487 95 496 97
rect 498 95 503 106
rect 505 101 510 106
rect 565 103 570 106
rect 563 102 570 103
rect 505 100 512 101
rect 505 96 507 100
rect 511 96 512 100
rect 563 98 564 102
rect 568 98 570 102
rect 563 97 570 98
rect 572 97 583 106
rect 505 95 512 96
rect 394 86 395 90
rect 399 86 401 90
rect 394 85 401 86
rect 487 90 494 95
rect 574 95 583 97
rect 585 95 590 106
rect 592 101 597 106
rect 1762 134 1772 136
rect 1762 131 1766 134
rect 1765 130 1766 131
rect 1770 133 1772 134
rect 2047 145 2054 146
rect 2047 141 2048 145
rect 2052 141 2054 145
rect 2047 140 2054 141
rect 2056 145 2064 146
rect 2056 141 2058 145
rect 2062 141 2064 145
rect 2056 140 2064 141
rect 2066 145 2074 146
rect 2066 141 2068 145
rect 2072 141 2074 145
rect 2066 140 2074 141
rect 2076 145 2083 146
rect 2076 141 2078 145
rect 2082 141 2083 145
rect 2376 143 2377 147
rect 2381 143 2383 147
rect 2376 142 2383 143
rect 2385 147 2393 148
rect 2385 143 2387 147
rect 2391 143 2393 147
rect 2385 142 2393 143
rect 2395 147 2403 148
rect 2395 143 2397 147
rect 2401 143 2403 147
rect 2395 142 2403 143
rect 2405 147 2412 148
rect 2405 143 2407 147
rect 2411 143 2412 147
rect 2703 146 2704 150
rect 2708 146 2710 150
rect 2703 145 2710 146
rect 2712 150 2720 151
rect 2712 146 2714 150
rect 2718 146 2720 150
rect 2712 145 2720 146
rect 2722 150 2730 151
rect 2722 146 2724 150
rect 2728 146 2730 150
rect 2722 145 2730 146
rect 2732 150 2739 151
rect 2732 146 2734 150
rect 2738 146 2739 150
rect 2732 145 2739 146
rect 2405 142 2412 143
rect 2076 140 2083 141
rect 1770 130 1779 133
rect 1765 128 1779 130
rect 1765 124 1779 126
rect 1765 120 1774 124
rect 1778 120 1779 124
rect 1765 118 1779 120
rect 1765 114 1779 116
rect 1765 110 1767 114
rect 1771 110 1774 114
rect 1778 110 1779 114
rect 1765 109 1779 110
rect 592 100 599 101
rect 592 96 594 100
rect 598 96 599 100
rect 592 95 599 96
rect 487 86 488 90
rect 492 86 494 90
rect 487 85 494 86
rect 574 90 581 95
rect 1738 108 1744 109
rect 1738 104 1739 108
rect 1743 107 1744 108
rect 1743 104 1747 107
rect 1738 102 1747 104
rect 1766 104 1772 105
rect 1766 103 1767 104
rect 1759 100 1767 103
rect 1771 103 1772 104
rect 1771 100 1779 103
rect 1738 95 1747 100
rect 1759 98 1779 100
rect 1738 91 1747 93
rect 1759 91 1779 96
rect 574 86 575 90
rect 579 86 581 90
rect 574 85 581 86
rect 1735 90 1753 91
rect 1735 86 1748 90
rect 1752 86 1753 90
rect 1735 85 1753 86
rect 1759 87 1779 89
rect 1735 83 1741 85
rect 1759 83 1760 87
rect 1764 83 1779 87
rect 1759 82 1779 83
rect 1735 79 1741 81
rect 1735 75 1736 79
rect 1740 75 1741 79
rect 1759 80 1773 82
rect 1759 76 1773 78
rect 1735 74 1741 75
rect 1759 73 1767 76
rect 1766 72 1767 73
rect 1771 72 1773 76
rect 1766 71 1773 72
rect 2250 32 2255 35
rect 2248 31 2255 32
rect 2248 27 2249 31
rect 2253 27 2255 31
rect 2248 26 2255 27
rect 2257 26 2268 35
rect 2259 24 2268 26
rect 2270 24 2275 35
rect 2277 30 2282 35
rect 2343 32 2348 35
rect 2341 31 2348 32
rect 2277 29 2284 30
rect 2277 25 2279 29
rect 2283 25 2284 29
rect 2341 27 2342 31
rect 2346 27 2348 31
rect 2341 26 2348 27
rect 2350 26 2361 35
rect 2277 24 2284 25
rect 2259 19 2266 24
rect 2352 24 2361 26
rect 2363 24 2368 35
rect 2370 30 2375 35
rect 2430 32 2435 35
rect 2428 31 2435 32
rect 2370 29 2377 30
rect 2370 25 2372 29
rect 2376 25 2377 29
rect 2428 27 2429 31
rect 2433 27 2435 31
rect 2428 26 2435 27
rect 2437 26 2448 35
rect 2370 24 2377 25
rect 2259 15 2260 19
rect 2264 15 2266 19
rect 2259 14 2266 15
rect 2352 19 2359 24
rect 2439 24 2448 26
rect 2450 24 2455 35
rect 2457 30 2462 35
rect 2457 29 2464 30
rect 2457 25 2459 29
rect 2463 25 2464 29
rect 2457 24 2464 25
rect 2352 15 2353 19
rect 2357 15 2359 19
rect 2352 14 2359 15
rect 2439 19 2446 24
rect 2439 15 2440 19
rect 2444 15 2446 19
rect 2439 14 2446 15
<< pdiffusion >>
rect 1714 1057 1724 1058
rect 1714 1053 1715 1057
rect 1719 1053 1724 1057
rect 1714 1051 1724 1053
rect 1714 1047 1724 1049
rect 1714 1043 1719 1047
rect 1723 1043 1724 1047
rect 1714 1041 1724 1043
rect 1054 1017 1085 1018
rect 1054 1013 1059 1017
rect 1063 1013 1085 1017
rect 1054 1012 1085 1013
rect 1087 1013 1103 1018
rect 1648 1028 1654 1029
rect 1714 1037 1724 1039
rect 1712 1033 1719 1037
rect 1723 1033 1724 1037
rect 1712 1031 1724 1033
rect 1648 1024 1649 1028
rect 1653 1027 1654 1028
rect 1653 1024 1660 1027
rect 1648 1022 1660 1024
rect 1712 1027 1724 1029
rect 1712 1024 1719 1027
rect 1718 1023 1719 1024
rect 1723 1023 1724 1027
rect 1109 1013 1122 1018
rect 1087 1012 1122 1013
rect 1142 1017 1157 1018
rect 1146 1013 1157 1017
rect 1142 1012 1157 1013
rect 1159 1017 1179 1018
rect 1159 1013 1175 1017
rect 1159 1012 1179 1013
rect 1186 1017 1196 1018
rect 1186 1013 1188 1017
rect 1192 1013 1196 1017
rect 1186 1012 1196 1013
rect 1198 1017 1217 1018
rect 1198 1013 1205 1017
rect 1209 1013 1217 1017
rect 1198 1012 1217 1013
rect 1219 1017 1227 1018
rect 1219 1013 1222 1017
rect 1226 1013 1227 1017
rect 1219 1012 1227 1013
rect 1240 1017 1250 1018
rect 1240 1013 1242 1017
rect 1246 1013 1250 1017
rect 1240 1012 1250 1013
rect 1252 1017 1271 1018
rect 1252 1013 1259 1017
rect 1263 1013 1271 1017
rect 1252 1012 1271 1013
rect 1273 1017 1281 1018
rect 1273 1013 1276 1017
rect 1280 1013 1281 1017
rect 1273 1012 1281 1013
rect 1296 1017 1306 1018
rect 1296 1013 1298 1017
rect 1302 1013 1306 1017
rect 1296 1012 1306 1013
rect 1308 1017 1327 1018
rect 1308 1013 1315 1017
rect 1319 1013 1327 1017
rect 1308 1012 1327 1013
rect 1329 1017 1337 1018
rect 1329 1013 1332 1017
rect 1336 1013 1337 1017
rect 1329 1012 1337 1013
rect 1350 1017 1360 1018
rect 1350 1013 1352 1017
rect 1356 1013 1360 1017
rect 1350 1012 1360 1013
rect 1362 1017 1381 1018
rect 1362 1013 1369 1017
rect 1373 1013 1381 1017
rect 1362 1012 1381 1013
rect 1383 1017 1391 1018
rect 1383 1013 1386 1017
rect 1390 1013 1391 1017
rect 1383 1012 1391 1013
rect 1648 1018 1660 1020
rect 1648 1014 1649 1018
rect 1653 1014 1660 1018
rect 1648 1012 1658 1014
rect 1718 1022 1724 1023
rect 178 987 184 994
rect 157 979 164 987
rect 157 975 158 979
rect 162 975 164 979
rect 157 974 164 975
rect 166 986 174 987
rect 166 982 168 986
rect 172 982 174 986
rect 166 979 174 982
rect 166 975 168 979
rect 172 975 174 979
rect 166 974 174 975
rect 176 981 184 987
rect 176 977 178 981
rect 182 977 184 981
rect 176 976 184 977
rect 186 993 193 994
rect 186 989 188 993
rect 192 989 193 993
rect 186 986 193 989
rect 265 987 271 994
rect 186 982 188 986
rect 192 982 193 986
rect 186 981 193 982
rect 186 976 191 981
rect 244 979 251 987
rect 176 974 182 976
rect 244 975 245 979
rect 249 975 251 979
rect 244 974 251 975
rect 253 986 261 987
rect 253 982 255 986
rect 259 982 261 986
rect 253 979 261 982
rect 253 975 255 979
rect 259 975 261 979
rect 253 974 261 975
rect 263 981 271 987
rect 263 977 265 981
rect 269 977 271 981
rect 263 976 271 977
rect 273 993 280 994
rect 273 989 275 993
rect 279 989 280 993
rect 273 986 280 989
rect 577 995 584 996
rect 358 987 364 994
rect 273 982 275 986
rect 279 982 280 986
rect 273 981 280 982
rect 273 976 278 981
rect 337 979 344 987
rect 263 974 269 976
rect 337 975 338 979
rect 342 975 344 979
rect 337 974 344 975
rect 346 986 354 987
rect 346 982 348 986
rect 352 982 354 986
rect 346 979 354 982
rect 346 975 348 979
rect 352 975 354 979
rect 346 974 354 975
rect 356 981 364 987
rect 356 977 358 981
rect 362 977 364 981
rect 356 976 364 977
rect 366 993 373 994
rect 366 989 368 993
rect 372 989 373 993
rect 366 986 373 989
rect 366 982 368 986
rect 372 982 373 986
rect 577 991 578 995
rect 582 991 584 995
rect 577 988 584 991
rect 577 984 578 988
rect 582 984 584 988
rect 577 983 584 984
rect 366 981 373 982
rect 366 976 371 981
rect 579 978 584 983
rect 586 989 592 996
rect 670 995 677 996
rect 670 991 671 995
rect 675 991 677 995
rect 586 983 594 989
rect 586 979 588 983
rect 592 979 594 983
rect 586 978 594 979
rect 356 974 362 976
rect 588 976 594 978
rect 596 988 604 989
rect 596 984 598 988
rect 602 984 604 988
rect 596 981 604 984
rect 596 977 598 981
rect 602 977 604 981
rect 596 976 604 977
rect 606 981 613 989
rect 670 988 677 991
rect 670 984 671 988
rect 675 984 677 988
rect 670 983 677 984
rect 606 977 608 981
rect 612 977 613 981
rect 672 978 677 983
rect 679 989 685 996
rect 757 995 764 996
rect 757 991 758 995
rect 762 991 764 995
rect 679 983 687 989
rect 679 979 681 983
rect 685 979 687 983
rect 679 978 687 979
rect 606 976 613 977
rect 681 976 687 978
rect 689 988 697 989
rect 689 984 691 988
rect 695 984 697 988
rect 689 981 697 984
rect 689 977 691 981
rect 695 977 697 981
rect 689 976 697 977
rect 699 981 706 989
rect 757 988 764 991
rect 757 984 758 988
rect 762 984 764 988
rect 757 983 764 984
rect 699 977 701 981
rect 705 977 706 981
rect 759 978 764 983
rect 766 989 772 996
rect 1648 1008 1658 1010
rect 1648 1004 1649 1008
rect 1653 1004 1658 1008
rect 1702 1011 1708 1012
rect 1702 1010 1703 1011
rect 1648 1002 1658 1004
rect 766 983 774 989
rect 766 979 768 983
rect 772 979 774 983
rect 766 978 774 979
rect 699 976 706 977
rect 768 976 774 978
rect 776 988 784 989
rect 776 984 778 988
rect 782 984 784 988
rect 776 981 784 984
rect 776 977 778 981
rect 782 977 784 981
rect 776 976 784 977
rect 786 981 793 989
rect 786 977 788 981
rect 792 977 793 981
rect 786 976 793 977
rect 1648 998 1658 1000
rect 1648 994 1653 998
rect 1657 994 1658 998
rect 1696 1007 1703 1010
rect 1707 1010 1708 1011
rect 1707 1007 1723 1010
rect 1696 1005 1723 1007
rect 1696 1001 1723 1003
rect 1696 998 1711 1001
rect 1705 997 1711 998
rect 1715 997 1723 1001
rect 1705 995 1723 997
rect 1648 993 1658 994
rect 1705 991 1723 993
rect 1705 987 1718 991
rect 1722 987 1723 991
rect 1705 985 1723 987
rect 1705 981 1723 983
rect 1696 975 1723 981
rect 1696 971 1697 975
rect 1701 971 1704 975
rect 1708 971 1723 975
rect 1696 969 1723 971
rect 1696 965 1723 967
rect 1696 962 1718 965
rect 1717 961 1718 962
rect 1722 961 1723 965
rect 1717 960 1723 961
rect 81 926 86 932
rect 79 925 86 926
rect 79 921 80 925
rect 84 921 86 925
rect 79 920 86 921
rect 88 930 94 932
rect 88 925 96 930
rect 88 921 90 925
rect 94 921 96 925
rect 88 920 96 921
rect 98 925 106 930
rect 98 921 100 925
rect 104 921 106 925
rect 98 920 106 921
rect 108 929 115 930
rect 108 925 110 929
rect 114 925 115 929
rect 167 927 172 948
rect 108 920 115 925
rect 165 926 172 927
rect 165 922 166 926
rect 170 922 172 926
rect 165 921 172 922
rect 174 947 186 948
rect 174 943 176 947
rect 180 943 186 947
rect 174 940 186 943
rect 174 936 176 940
rect 180 939 186 940
rect 203 939 208 948
rect 180 936 188 939
rect 174 921 188 936
rect 190 926 198 939
rect 190 922 192 926
rect 196 922 198 926
rect 190 921 198 922
rect 200 933 208 939
rect 200 929 202 933
rect 206 929 208 933
rect 200 921 208 929
rect 210 942 215 948
rect 210 941 217 942
rect 210 937 212 941
rect 216 937 217 941
rect 210 936 217 937
rect 210 921 215 936
rect 251 927 256 948
rect 249 926 256 927
rect 249 922 250 926
rect 254 922 256 926
rect 249 921 256 922
rect 258 947 270 948
rect 258 943 260 947
rect 264 943 270 947
rect 258 940 270 943
rect 258 936 260 940
rect 264 939 270 940
rect 287 939 292 948
rect 264 936 272 939
rect 258 921 272 936
rect 274 926 282 939
rect 274 922 276 926
rect 280 922 282 926
rect 274 921 282 922
rect 284 933 292 939
rect 284 929 286 933
rect 290 929 292 933
rect 284 921 292 929
rect 294 942 299 948
rect 294 941 301 942
rect 294 937 296 941
rect 300 937 301 941
rect 294 936 301 937
rect 294 921 299 936
rect 313 926 318 932
rect 311 925 318 926
rect 311 921 312 925
rect 316 921 318 925
rect 311 920 318 921
rect 320 930 326 932
rect 320 925 328 930
rect 320 921 322 925
rect 326 921 328 925
rect 320 920 328 921
rect 330 925 338 930
rect 330 921 332 925
rect 336 921 338 925
rect 330 920 338 921
rect 340 929 347 930
rect 340 925 342 929
rect 346 925 347 929
rect 410 928 415 934
rect 340 920 347 925
rect 408 927 415 928
rect 408 923 409 927
rect 413 923 415 927
rect 408 922 415 923
rect 417 932 423 934
rect 417 927 425 932
rect 417 923 419 927
rect 423 923 425 927
rect 417 922 425 923
rect 427 927 435 932
rect 427 923 429 927
rect 433 923 435 927
rect 427 922 435 923
rect 437 931 444 932
rect 437 927 439 931
rect 443 927 444 931
rect 496 929 501 950
rect 437 922 444 927
rect 494 928 501 929
rect 494 924 495 928
rect 499 924 501 928
rect 494 923 501 924
rect 503 949 515 950
rect 503 945 505 949
rect 509 945 515 949
rect 503 942 515 945
rect 503 938 505 942
rect 509 941 515 942
rect 532 941 537 950
rect 509 938 517 941
rect 503 923 517 938
rect 519 928 527 941
rect 519 924 521 928
rect 525 924 527 928
rect 519 923 527 924
rect 529 935 537 941
rect 529 931 531 935
rect 535 931 537 935
rect 529 923 537 931
rect 539 944 544 950
rect 539 943 546 944
rect 539 939 541 943
rect 545 939 546 943
rect 539 938 546 939
rect 539 923 544 938
rect 580 929 585 950
rect 578 928 585 929
rect 578 924 579 928
rect 583 924 585 928
rect 578 923 585 924
rect 587 949 599 950
rect 587 945 589 949
rect 593 945 599 949
rect 587 942 599 945
rect 587 938 589 942
rect 593 941 599 942
rect 616 941 621 950
rect 593 938 601 941
rect 587 923 601 938
rect 603 928 611 941
rect 603 924 605 928
rect 609 924 611 928
rect 603 923 611 924
rect 613 935 621 941
rect 613 931 615 935
rect 619 931 621 935
rect 613 923 621 931
rect 623 944 628 950
rect 623 943 630 944
rect 623 939 625 943
rect 629 939 630 943
rect 623 938 630 939
rect 623 923 628 938
rect 642 928 647 934
rect 640 927 647 928
rect 640 923 641 927
rect 645 923 647 927
rect 640 922 647 923
rect 649 932 655 934
rect 649 927 657 932
rect 649 923 651 927
rect 655 923 657 927
rect 649 922 657 923
rect 659 927 667 932
rect 659 923 661 927
rect 665 923 667 927
rect 659 922 667 923
rect 669 931 676 932
rect 737 931 742 937
rect 669 927 671 931
rect 675 927 676 931
rect 669 922 676 927
rect 735 930 742 931
rect 735 926 736 930
rect 740 926 742 930
rect 735 925 742 926
rect 744 935 750 937
rect 744 930 752 935
rect 744 926 746 930
rect 750 926 752 930
rect 744 925 752 926
rect 754 930 762 935
rect 754 926 756 930
rect 760 926 762 930
rect 754 925 762 926
rect 764 934 771 935
rect 764 930 766 934
rect 770 930 771 934
rect 823 932 828 953
rect 764 925 771 930
rect 821 931 828 932
rect 821 927 822 931
rect 826 927 828 931
rect 821 926 828 927
rect 830 952 842 953
rect 830 948 832 952
rect 836 948 842 952
rect 830 945 842 948
rect 830 941 832 945
rect 836 944 842 945
rect 859 944 864 953
rect 836 941 844 944
rect 830 926 844 941
rect 846 931 854 944
rect 846 927 848 931
rect 852 927 854 931
rect 846 926 854 927
rect 856 938 864 944
rect 856 934 858 938
rect 862 934 864 938
rect 856 926 864 934
rect 866 947 871 953
rect 866 946 873 947
rect 866 942 868 946
rect 872 942 873 946
rect 866 941 873 942
rect 866 926 871 941
rect 907 932 912 953
rect 905 931 912 932
rect 905 927 906 931
rect 910 927 912 931
rect 905 926 912 927
rect 914 952 926 953
rect 914 948 916 952
rect 920 948 926 952
rect 914 945 926 948
rect 914 941 916 945
rect 920 944 926 945
rect 943 944 948 953
rect 920 941 928 944
rect 914 926 928 941
rect 930 931 938 944
rect 930 927 932 931
rect 936 927 938 931
rect 930 926 938 927
rect 940 938 948 944
rect 940 934 942 938
rect 946 934 948 938
rect 940 926 948 934
rect 950 947 955 953
rect 950 946 957 947
rect 950 942 952 946
rect 956 942 957 946
rect 950 941 957 942
rect 950 926 955 941
rect 969 931 974 937
rect 967 930 974 931
rect 967 926 968 930
rect 972 926 974 930
rect 967 925 974 926
rect 976 935 982 937
rect 976 930 984 935
rect 976 926 978 930
rect 982 926 984 930
rect 976 925 984 926
rect 986 930 994 935
rect 986 926 988 930
rect 992 926 994 930
rect 986 925 994 926
rect 996 934 1003 935
rect 996 930 998 934
rect 1002 930 1003 934
rect 1553 935 1559 936
rect 1553 934 1554 935
rect 996 925 1003 930
rect 1546 931 1554 934
rect 1558 934 1559 935
rect 1558 931 1564 934
rect 1546 929 1564 931
rect 1546 922 1564 927
rect 1146 918 1161 919
rect 1150 914 1161 918
rect 1146 913 1161 914
rect 1163 918 1183 919
rect 1163 914 1179 918
rect 1163 913 1183 914
rect 1190 918 1200 919
rect 1190 914 1192 918
rect 1196 914 1200 918
rect 1190 913 1200 914
rect 1202 918 1221 919
rect 1202 914 1209 918
rect 1213 914 1221 918
rect 1202 913 1221 914
rect 1223 918 1231 919
rect 1223 914 1226 918
rect 1230 914 1231 918
rect 1223 913 1231 914
rect 1244 918 1254 919
rect 1244 914 1246 918
rect 1250 914 1254 918
rect 1244 913 1254 914
rect 1256 918 1275 919
rect 1256 914 1263 918
rect 1267 914 1275 918
rect 1256 913 1275 914
rect 1277 918 1285 919
rect 1277 914 1280 918
rect 1284 914 1285 918
rect 1277 913 1285 914
rect 1300 918 1310 919
rect 1300 914 1302 918
rect 1306 914 1310 918
rect 1300 913 1310 914
rect 1312 918 1331 919
rect 1312 914 1319 918
rect 1323 914 1331 918
rect 1312 913 1331 914
rect 1333 918 1341 919
rect 1333 914 1336 918
rect 1340 914 1341 918
rect 1333 913 1341 914
rect 1354 918 1364 919
rect 1354 914 1356 918
rect 1360 914 1364 918
rect 1354 913 1364 914
rect 1366 918 1385 919
rect 1366 914 1373 918
rect 1377 914 1385 918
rect 1366 913 1385 914
rect 1387 918 1395 919
rect 1387 914 1390 918
rect 1394 914 1395 918
rect 1387 913 1395 914
rect 1546 917 1564 920
rect 1546 913 1547 917
rect 1551 913 1567 917
rect 1546 911 1567 913
rect 1555 909 1567 911
rect 1555 905 1567 907
rect 1555 901 1556 905
rect 1560 902 1567 905
rect 1560 901 1561 902
rect 1555 900 1561 901
rect 1649 942 1655 943
rect 1649 938 1650 942
rect 1654 941 1655 942
rect 1654 938 1676 941
rect 1649 936 1676 938
rect 1649 932 1676 934
rect 1649 928 1664 932
rect 1668 928 1671 932
rect 1675 928 1676 932
rect 1649 922 1676 928
rect 1702 927 1708 928
rect 1702 926 1703 927
rect 1696 923 1703 926
rect 1707 926 1708 927
rect 1707 923 1723 926
rect 1649 920 1667 922
rect 1696 921 1723 923
rect 2462 927 2471 928
rect 2462 923 2464 927
rect 2468 923 2471 927
rect 1649 916 1667 918
rect 1696 917 1723 919
rect 1649 912 1650 916
rect 1654 912 1667 916
rect 1649 910 1667 912
rect 1696 914 1711 917
rect 1705 913 1711 914
rect 1715 913 1723 917
rect 2462 919 2471 923
rect 1705 911 1723 913
rect 1649 906 1667 908
rect 1649 902 1657 906
rect 1661 905 1667 906
rect 1661 902 1676 905
rect 1705 907 1723 909
rect 1705 903 1718 907
rect 1722 903 1723 907
rect 1649 900 1676 902
rect 1705 901 1723 903
rect 1649 896 1676 898
rect 1705 897 1723 899
rect 1649 893 1665 896
rect 1430 890 1436 891
rect 1430 886 1431 890
rect 1435 888 1436 890
rect 1664 892 1665 893
rect 1669 893 1676 896
rect 1669 892 1670 893
rect 1664 891 1670 892
rect 1696 891 1723 897
rect 1435 886 1438 888
rect 1054 872 1085 873
rect 1054 868 1059 872
rect 1063 868 1085 872
rect 191 836 199 839
rect 174 831 179 836
rect 172 830 179 831
rect 172 826 173 830
rect 177 826 179 830
rect 172 825 179 826
rect 174 818 179 825
rect 181 818 186 836
rect 188 827 199 836
rect 201 833 206 839
rect 1054 867 1085 868
rect 1087 868 1103 873
rect 1430 877 1438 886
rect 1421 873 1426 877
rect 1109 868 1122 873
rect 1087 867 1122 868
rect 1142 872 1157 873
rect 1146 868 1157 872
rect 1142 867 1157 868
rect 1159 872 1179 873
rect 1159 868 1175 872
rect 1159 867 1179 868
rect 1186 872 1196 873
rect 1186 868 1188 872
rect 1192 868 1196 872
rect 1186 867 1196 868
rect 1198 872 1217 873
rect 1198 868 1205 872
rect 1209 868 1217 872
rect 1198 867 1217 868
rect 1219 872 1227 873
rect 1219 868 1222 872
rect 1226 868 1227 872
rect 1219 867 1227 868
rect 1240 872 1250 873
rect 1240 868 1242 872
rect 1246 868 1250 872
rect 1240 867 1250 868
rect 1252 872 1271 873
rect 1252 868 1259 872
rect 1263 868 1271 872
rect 1252 867 1271 868
rect 1273 872 1281 873
rect 1273 868 1276 872
rect 1280 868 1281 872
rect 1273 867 1281 868
rect 1296 872 1306 873
rect 1296 868 1298 872
rect 1302 868 1306 872
rect 1296 867 1306 868
rect 1308 872 1327 873
rect 1308 868 1315 872
rect 1319 868 1327 872
rect 1308 867 1327 868
rect 1329 872 1337 873
rect 1329 868 1332 872
rect 1336 868 1337 872
rect 1329 867 1337 868
rect 1350 872 1360 873
rect 1350 868 1352 872
rect 1356 868 1360 872
rect 1350 867 1360 868
rect 1362 872 1381 873
rect 1362 868 1369 872
rect 1373 868 1381 872
rect 1362 867 1381 868
rect 1383 872 1391 873
rect 1383 868 1386 872
rect 1390 868 1391 872
rect 1383 867 1391 868
rect 1419 872 1426 873
rect 1419 868 1420 872
rect 1424 868 1426 872
rect 1419 867 1426 868
rect 1421 860 1426 867
rect 1428 860 1438 877
rect 1440 881 1445 888
rect 1696 887 1697 891
rect 1701 887 1704 891
rect 1708 887 1723 891
rect 1696 885 1723 887
rect 1696 881 1723 883
rect 1440 880 1447 881
rect 1440 876 1442 880
rect 1446 876 1447 880
rect 1696 878 1718 881
rect 1717 877 1718 878
rect 1722 877 1723 881
rect 1717 876 1723 877
rect 1811 918 1817 919
rect 2451 918 2458 919
rect 1811 917 1812 918
rect 1805 914 1812 917
rect 1816 914 1817 918
rect 1805 912 1817 914
rect 2451 914 2452 918
rect 2456 914 2458 918
rect 2451 913 2458 914
rect 1805 908 1817 910
rect 1805 906 1826 908
rect 2453 907 2458 913
rect 2460 910 2471 919
rect 2473 910 2478 928
rect 2480 921 2485 928
rect 2480 920 2487 921
rect 2480 916 2482 920
rect 2486 916 2487 920
rect 2680 918 2685 930
rect 2480 915 2487 916
rect 2678 917 2685 918
rect 2480 910 2485 915
rect 2678 913 2679 917
rect 2683 913 2685 917
rect 2678 910 2685 913
rect 2460 907 2468 910
rect 1805 902 1821 906
rect 1825 902 1826 906
rect 1808 899 1826 902
rect 1808 892 1826 897
rect 2678 906 2679 910
rect 2683 906 2685 910
rect 2678 905 2685 906
rect 2687 929 2696 930
rect 2687 925 2690 929
rect 2694 925 2696 929
rect 2719 929 2733 930
rect 2719 927 2725 929
rect 2687 918 2696 925
rect 2703 918 2708 927
rect 2687 905 2698 918
rect 2700 910 2708 918
rect 2700 906 2702 910
rect 2706 906 2708 910
rect 2700 905 2708 906
rect 1808 888 1826 890
rect 1808 885 1814 888
rect 1813 884 1814 885
rect 1818 885 1826 888
rect 1818 884 1819 885
rect 1813 883 1819 884
rect 2703 902 2708 905
rect 2710 902 2715 927
rect 2717 925 2725 927
rect 2729 925 2733 929
rect 2717 922 2733 925
rect 2717 918 2725 922
rect 2729 918 2733 922
rect 2717 902 2733 918
rect 2735 921 2743 930
rect 2735 917 2737 921
rect 2741 917 2743 921
rect 2735 914 2743 917
rect 2735 910 2737 914
rect 2741 910 2743 914
rect 2735 902 2743 910
rect 2745 929 2753 930
rect 2745 925 2747 929
rect 2751 925 2753 929
rect 2745 922 2753 925
rect 2745 918 2747 922
rect 2751 918 2753 922
rect 2745 902 2753 918
rect 2755 915 2760 930
rect 2822 929 2831 930
rect 2822 925 2824 929
rect 2828 925 2831 929
rect 2822 921 2831 925
rect 2811 920 2818 921
rect 2811 916 2812 920
rect 2816 916 2818 920
rect 2811 915 2818 916
rect 2755 914 2762 915
rect 2755 910 2757 914
rect 2761 910 2762 914
rect 2755 907 2762 910
rect 2813 909 2818 915
rect 2820 912 2831 921
rect 2833 912 2838 930
rect 2840 923 2845 930
rect 2840 922 2847 923
rect 2840 918 2842 922
rect 2846 918 2847 922
rect 2840 917 2847 918
rect 2840 912 2845 917
rect 2820 909 2828 912
rect 2755 903 2757 907
rect 2761 903 2762 907
rect 2755 902 2762 903
rect 1440 873 1447 876
rect 1440 869 1442 873
rect 1446 869 1447 873
rect 1440 868 1447 869
rect 1440 860 1445 868
rect 847 841 855 844
rect 520 838 528 841
rect 503 833 508 838
rect 201 832 208 833
rect 201 828 203 832
rect 207 828 208 832
rect 201 827 208 828
rect 501 832 508 833
rect 501 828 502 832
rect 506 828 508 832
rect 501 827 508 828
rect 188 823 197 827
rect 188 819 191 823
rect 195 819 197 823
rect 188 818 197 819
rect 503 820 508 827
rect 510 820 515 838
rect 517 829 528 838
rect 530 835 535 841
rect 830 836 835 841
rect 828 835 835 836
rect 530 834 537 835
rect 530 830 532 834
rect 536 830 537 834
rect 828 831 829 835
rect 833 831 835 835
rect 828 830 835 831
rect 530 829 537 830
rect 517 825 526 829
rect 517 821 520 825
rect 524 821 526 825
rect 830 823 835 830
rect 837 823 842 841
rect 844 832 855 841
rect 857 838 862 844
rect 857 837 864 838
rect 857 833 859 837
rect 863 833 864 837
rect 857 832 864 833
rect 844 828 853 832
rect 1649 858 1655 859
rect 1649 854 1650 858
rect 1654 857 1655 858
rect 1654 854 1676 857
rect 1649 852 1676 854
rect 1649 848 1676 850
rect 1649 844 1664 848
rect 1668 844 1671 848
rect 1675 844 1676 848
rect 1649 838 1676 844
rect 1649 836 1667 838
rect 844 824 847 828
rect 851 824 853 828
rect 1649 832 1667 834
rect 844 823 853 824
rect 517 820 526 821
rect 1649 828 1650 832
rect 1654 828 1667 832
rect 1649 826 1667 828
rect 1714 825 1724 826
rect 1649 822 1667 824
rect 80 780 85 786
rect 78 779 85 780
rect 78 775 79 779
rect 83 775 85 779
rect 78 774 85 775
rect 87 784 93 786
rect 87 779 95 784
rect 87 775 89 779
rect 93 775 95 779
rect 87 774 95 775
rect 97 779 105 784
rect 97 775 99 779
rect 103 775 105 779
rect 97 774 105 775
rect 107 783 114 784
rect 107 779 109 783
rect 113 779 114 783
rect 166 781 171 802
rect 107 774 114 779
rect 164 780 171 781
rect 164 776 165 780
rect 169 776 171 780
rect 164 775 171 776
rect 173 801 185 802
rect 173 797 175 801
rect 179 797 185 801
rect 173 794 185 797
rect 173 790 175 794
rect 179 793 185 794
rect 202 793 207 802
rect 179 790 187 793
rect 173 775 187 790
rect 189 780 197 793
rect 189 776 191 780
rect 195 776 197 780
rect 189 775 197 776
rect 199 787 207 793
rect 199 783 201 787
rect 205 783 207 787
rect 199 775 207 783
rect 209 796 214 802
rect 209 795 216 796
rect 209 791 211 795
rect 215 791 216 795
rect 209 790 216 791
rect 209 775 214 790
rect 250 781 255 802
rect 248 780 255 781
rect 248 776 249 780
rect 253 776 255 780
rect 248 775 255 776
rect 257 801 269 802
rect 257 797 259 801
rect 263 797 269 801
rect 257 794 269 797
rect 257 790 259 794
rect 263 793 269 794
rect 286 793 291 802
rect 263 790 271 793
rect 257 775 271 790
rect 273 780 281 793
rect 273 776 275 780
rect 279 776 281 780
rect 273 775 281 776
rect 283 787 291 793
rect 283 783 285 787
rect 289 783 291 787
rect 283 775 291 783
rect 293 796 298 802
rect 293 795 300 796
rect 293 791 295 795
rect 299 791 300 795
rect 293 790 300 791
rect 293 775 298 790
rect 312 780 317 786
rect 310 779 317 780
rect 310 775 311 779
rect 315 775 317 779
rect 310 774 317 775
rect 319 784 325 786
rect 319 779 327 784
rect 319 775 321 779
rect 325 775 327 779
rect 319 774 327 775
rect 329 779 337 784
rect 329 775 331 779
rect 335 775 337 779
rect 329 774 337 775
rect 339 783 346 784
rect 339 779 341 783
rect 345 779 346 783
rect 409 782 414 788
rect 339 774 346 779
rect 407 781 414 782
rect 407 777 408 781
rect 412 777 414 781
rect 407 776 414 777
rect 416 786 422 788
rect 416 781 424 786
rect 416 777 418 781
rect 422 777 424 781
rect 416 776 424 777
rect 426 781 434 786
rect 426 777 428 781
rect 432 777 434 781
rect 426 776 434 777
rect 436 785 443 786
rect 436 781 438 785
rect 442 781 443 785
rect 495 783 500 804
rect 436 776 443 781
rect 493 782 500 783
rect 493 778 494 782
rect 498 778 500 782
rect 493 777 500 778
rect 502 803 514 804
rect 502 799 504 803
rect 508 799 514 803
rect 502 796 514 799
rect 502 792 504 796
rect 508 795 514 796
rect 531 795 536 804
rect 508 792 516 795
rect 502 777 516 792
rect 518 782 526 795
rect 518 778 520 782
rect 524 778 526 782
rect 518 777 526 778
rect 528 789 536 795
rect 528 785 530 789
rect 534 785 536 789
rect 528 777 536 785
rect 538 798 543 804
rect 538 797 545 798
rect 538 793 540 797
rect 544 793 545 797
rect 538 792 545 793
rect 538 777 543 792
rect 579 783 584 804
rect 577 782 584 783
rect 577 778 578 782
rect 582 778 584 782
rect 577 777 584 778
rect 586 803 598 804
rect 586 799 588 803
rect 592 799 598 803
rect 586 796 598 799
rect 586 792 588 796
rect 592 795 598 796
rect 615 795 620 804
rect 592 792 600 795
rect 586 777 600 792
rect 602 782 610 795
rect 602 778 604 782
rect 608 778 610 782
rect 602 777 610 778
rect 612 789 620 795
rect 612 785 614 789
rect 618 785 620 789
rect 612 777 620 785
rect 622 798 627 804
rect 622 797 629 798
rect 622 793 624 797
rect 628 793 629 797
rect 622 792 629 793
rect 622 777 627 792
rect 641 782 646 788
rect 639 781 646 782
rect 639 777 640 781
rect 644 777 646 781
rect 639 776 646 777
rect 648 786 654 788
rect 648 781 656 786
rect 648 777 650 781
rect 654 777 656 781
rect 648 776 656 777
rect 658 781 666 786
rect 658 777 660 781
rect 664 777 666 781
rect 658 776 666 777
rect 668 785 675 786
rect 736 785 741 791
rect 668 781 670 785
rect 674 781 675 785
rect 668 776 675 781
rect 734 784 741 785
rect 734 780 735 784
rect 739 780 741 784
rect 734 779 741 780
rect 743 789 749 791
rect 743 784 751 789
rect 743 780 745 784
rect 749 780 751 784
rect 743 779 751 780
rect 753 784 761 789
rect 753 780 755 784
rect 759 780 761 784
rect 753 779 761 780
rect 763 788 770 789
rect 763 784 765 788
rect 769 784 770 788
rect 822 786 827 807
rect 763 779 770 784
rect 820 785 827 786
rect 820 781 821 785
rect 825 781 827 785
rect 820 780 827 781
rect 829 806 841 807
rect 829 802 831 806
rect 835 802 841 806
rect 829 799 841 802
rect 829 795 831 799
rect 835 798 841 799
rect 858 798 863 807
rect 835 795 843 798
rect 829 780 843 795
rect 845 785 853 798
rect 845 781 847 785
rect 851 781 853 785
rect 845 780 853 781
rect 855 792 863 798
rect 855 788 857 792
rect 861 788 863 792
rect 855 780 863 788
rect 865 801 870 807
rect 865 800 872 801
rect 865 796 867 800
rect 871 796 872 800
rect 865 795 872 796
rect 865 780 870 795
rect 906 786 911 807
rect 904 785 911 786
rect 904 781 905 785
rect 909 781 911 785
rect 904 780 911 781
rect 913 806 925 807
rect 913 802 915 806
rect 919 802 925 806
rect 913 799 925 802
rect 913 795 915 799
rect 919 798 925 799
rect 942 798 947 807
rect 919 795 927 798
rect 913 780 927 795
rect 929 785 937 798
rect 929 781 931 785
rect 935 781 937 785
rect 929 780 937 781
rect 939 792 947 798
rect 939 788 941 792
rect 945 788 947 792
rect 939 780 947 788
rect 949 801 954 807
rect 949 800 956 801
rect 949 796 951 800
rect 955 796 956 800
rect 949 795 956 796
rect 949 780 954 795
rect 968 785 973 791
rect 966 784 973 785
rect 966 780 967 784
rect 971 780 973 784
rect 966 779 973 780
rect 975 789 981 791
rect 1649 818 1657 822
rect 1661 821 1667 822
rect 1661 818 1676 821
rect 1649 816 1676 818
rect 1649 812 1676 814
rect 1649 809 1665 812
rect 1664 808 1665 809
rect 1669 809 1676 812
rect 1714 821 1715 825
rect 1719 821 1724 825
rect 1714 819 1724 821
rect 2312 821 2319 826
rect 1714 815 1724 817
rect 2312 817 2313 821
rect 2317 817 2319 821
rect 2312 816 2319 817
rect 2321 825 2329 826
rect 2321 821 2323 825
rect 2327 821 2329 825
rect 2321 816 2329 821
rect 2331 825 2339 826
rect 2331 821 2333 825
rect 2337 821 2339 825
rect 2331 816 2339 821
rect 1669 808 1670 809
rect 1664 807 1670 808
rect 1714 811 1719 815
rect 1723 811 1724 815
rect 2333 814 2339 816
rect 2341 825 2348 826
rect 2341 821 2343 825
rect 2347 821 2348 825
rect 2341 820 2348 821
rect 2341 814 2346 820
rect 1714 809 1724 811
rect 1648 796 1654 797
rect 1714 805 1724 807
rect 1712 801 1719 805
rect 1723 801 1724 805
rect 1712 799 1724 801
rect 2360 810 2365 825
rect 2358 809 2365 810
rect 2358 805 2359 809
rect 2363 805 2365 809
rect 2358 804 2365 805
rect 1648 792 1649 796
rect 1653 795 1654 796
rect 1653 792 1660 795
rect 1648 790 1660 792
rect 1712 795 1724 797
rect 1712 792 1719 795
rect 1718 791 1719 792
rect 1723 791 1724 795
rect 975 784 983 789
rect 975 780 977 784
rect 981 780 983 784
rect 975 779 983 780
rect 985 784 993 789
rect 985 780 987 784
rect 991 780 993 784
rect 985 779 993 780
rect 995 788 1002 789
rect 995 784 997 788
rect 1001 784 1002 788
rect 995 779 1002 784
rect 1422 780 1427 787
rect 1420 779 1427 780
rect 1420 775 1421 779
rect 1425 775 1427 779
rect 1420 774 1427 775
rect 1146 773 1161 774
rect 1150 769 1161 773
rect 1146 768 1161 769
rect 1163 773 1183 774
rect 1163 769 1179 773
rect 1163 768 1183 769
rect 1190 773 1200 774
rect 1190 769 1192 773
rect 1196 769 1200 773
rect 1190 768 1200 769
rect 1202 773 1221 774
rect 1202 769 1209 773
rect 1213 769 1221 773
rect 1202 768 1221 769
rect 1223 773 1231 774
rect 1223 769 1226 773
rect 1230 769 1231 773
rect 1223 768 1231 769
rect 1244 773 1254 774
rect 1244 769 1246 773
rect 1250 769 1254 773
rect 1244 768 1254 769
rect 1256 773 1275 774
rect 1256 769 1263 773
rect 1267 769 1275 773
rect 1256 768 1275 769
rect 1277 773 1285 774
rect 1277 769 1280 773
rect 1284 769 1285 773
rect 1277 768 1285 769
rect 1300 773 1310 774
rect 1300 769 1302 773
rect 1306 769 1310 773
rect 1300 768 1310 769
rect 1312 773 1331 774
rect 1312 769 1319 773
rect 1323 769 1331 773
rect 1312 768 1331 769
rect 1333 773 1341 774
rect 1333 769 1336 773
rect 1340 769 1341 773
rect 1333 768 1341 769
rect 1354 773 1364 774
rect 1354 769 1356 773
rect 1360 769 1364 773
rect 1354 768 1364 769
rect 1366 773 1385 774
rect 1366 769 1373 773
rect 1377 769 1385 773
rect 1366 768 1385 769
rect 1387 773 1395 774
rect 1387 769 1390 773
rect 1394 769 1395 773
rect 1422 770 1427 774
rect 1429 770 1439 787
rect 1387 768 1395 769
rect 1431 761 1439 770
rect 1431 757 1432 761
rect 1436 759 1439 761
rect 1441 779 1446 787
rect 1648 786 1660 788
rect 1648 782 1649 786
rect 1653 782 1660 786
rect 1648 780 1658 782
rect 1718 790 1724 791
rect 2360 798 2365 804
rect 2367 817 2375 825
rect 2367 813 2369 817
rect 2373 813 2375 817
rect 2367 807 2375 813
rect 2377 824 2385 825
rect 2377 820 2379 824
rect 2383 820 2385 824
rect 2377 807 2385 820
rect 2387 810 2401 825
rect 2387 807 2395 810
rect 2367 798 2372 807
rect 2389 806 2395 807
rect 2399 806 2401 810
rect 2389 803 2401 806
rect 2389 799 2395 803
rect 2399 799 2401 803
rect 2389 798 2401 799
rect 2403 824 2410 825
rect 2403 820 2405 824
rect 2409 820 2410 824
rect 2403 819 2410 820
rect 2403 798 2408 819
rect 2444 810 2449 825
rect 2442 809 2449 810
rect 2442 805 2443 809
rect 2447 805 2449 809
rect 2442 804 2449 805
rect 2444 798 2449 804
rect 2451 817 2459 825
rect 2451 813 2453 817
rect 2457 813 2459 817
rect 2451 807 2459 813
rect 2461 824 2469 825
rect 2461 820 2463 824
rect 2467 820 2469 824
rect 2461 807 2469 820
rect 2471 810 2485 825
rect 2471 807 2479 810
rect 2451 798 2456 807
rect 2473 806 2479 807
rect 2483 806 2485 810
rect 2473 803 2485 806
rect 2473 799 2479 803
rect 2483 799 2485 803
rect 2473 798 2485 799
rect 2487 824 2494 825
rect 2487 820 2489 824
rect 2493 820 2494 824
rect 2487 819 2494 820
rect 2544 821 2551 826
rect 2487 798 2492 819
rect 2544 817 2545 821
rect 2549 817 2551 821
rect 2544 816 2551 817
rect 2553 825 2561 826
rect 2553 821 2555 825
rect 2559 821 2561 825
rect 2553 816 2561 821
rect 2563 825 2571 826
rect 2563 821 2565 825
rect 2569 821 2571 825
rect 2563 816 2571 821
rect 2565 814 2571 816
rect 2573 825 2580 826
rect 2573 821 2575 825
rect 2579 821 2580 825
rect 2573 820 2580 821
rect 2672 823 2679 828
rect 2573 814 2578 820
rect 2672 819 2673 823
rect 2677 819 2679 823
rect 2672 818 2679 819
rect 2681 827 2689 828
rect 2681 823 2683 827
rect 2687 823 2689 827
rect 2681 818 2689 823
rect 2691 827 2699 828
rect 2691 823 2693 827
rect 2697 823 2699 827
rect 2691 818 2699 823
rect 2693 816 2699 818
rect 2701 827 2708 828
rect 2701 823 2703 827
rect 2707 823 2708 827
rect 2701 822 2708 823
rect 2701 816 2706 822
rect 2720 812 2725 827
rect 2718 811 2725 812
rect 2718 807 2719 811
rect 2723 807 2725 811
rect 2718 806 2725 807
rect 2720 800 2725 806
rect 2727 819 2735 827
rect 2727 815 2729 819
rect 2733 815 2735 819
rect 2727 809 2735 815
rect 2737 826 2745 827
rect 2737 822 2739 826
rect 2743 822 2745 826
rect 2737 809 2745 822
rect 2747 812 2761 827
rect 2747 809 2755 812
rect 2727 800 2732 809
rect 2749 808 2755 809
rect 2759 808 2761 812
rect 2749 805 2761 808
rect 2749 801 2755 805
rect 2759 801 2761 805
rect 2749 800 2761 801
rect 2763 826 2770 827
rect 2763 822 2765 826
rect 2769 822 2770 826
rect 2763 821 2770 822
rect 2763 800 2768 821
rect 2804 812 2809 827
rect 2802 811 2809 812
rect 2802 807 2803 811
rect 2807 807 2809 811
rect 2802 806 2809 807
rect 2804 800 2809 806
rect 2811 819 2819 827
rect 2811 815 2813 819
rect 2817 815 2819 819
rect 2811 809 2819 815
rect 2821 826 2829 827
rect 2821 822 2823 826
rect 2827 822 2829 826
rect 2821 809 2829 822
rect 2831 812 2845 827
rect 2831 809 2839 812
rect 2811 800 2816 809
rect 2833 808 2839 809
rect 2843 808 2845 812
rect 2833 805 2845 808
rect 2833 801 2839 805
rect 2843 801 2845 805
rect 2833 800 2845 801
rect 2847 826 2854 827
rect 2847 822 2849 826
rect 2853 822 2854 826
rect 2847 821 2854 822
rect 2904 823 2911 828
rect 2847 800 2852 821
rect 2904 819 2905 823
rect 2909 819 2911 823
rect 2904 818 2911 819
rect 2913 827 2921 828
rect 2913 823 2915 827
rect 2919 823 2921 827
rect 2913 818 2921 823
rect 2923 827 2931 828
rect 2923 823 2925 827
rect 2929 823 2931 827
rect 2923 818 2931 823
rect 2925 816 2931 818
rect 2933 827 2940 828
rect 2933 823 2935 827
rect 2939 823 2940 827
rect 2933 822 2940 823
rect 2933 816 2938 822
rect 1441 778 1448 779
rect 1441 774 1443 778
rect 1447 774 1448 778
rect 1648 776 1658 778
rect 1441 771 1448 774
rect 1648 772 1649 776
rect 1653 772 1658 776
rect 1441 767 1443 771
rect 1447 767 1448 771
rect 1648 770 1658 772
rect 1441 766 1448 767
rect 1441 759 1446 766
rect 1648 766 1658 768
rect 1648 762 1653 766
rect 1657 762 1658 766
rect 1987 764 1992 770
rect 1985 763 1992 764
rect 1648 761 1658 762
rect 1985 759 1986 763
rect 1990 759 1992 763
rect 1436 757 1437 759
rect 1431 756 1437 757
rect 1985 758 1992 759
rect 1994 768 2000 770
rect 1994 763 2002 768
rect 1994 759 1996 763
rect 2000 759 2002 763
rect 1994 758 2002 759
rect 2004 763 2012 768
rect 2004 759 2006 763
rect 2010 759 2012 763
rect 2004 758 2012 759
rect 2014 767 2021 768
rect 2014 763 2016 767
rect 2020 763 2021 767
rect 2073 765 2078 786
rect 2014 758 2021 763
rect 1430 750 1436 751
rect 1430 746 1431 750
rect 1435 748 1436 750
rect 1435 746 1438 748
rect 1430 737 1438 746
rect 1053 730 1084 731
rect 1053 726 1058 730
rect 1062 726 1084 730
rect 1053 725 1084 726
rect 1086 726 1102 731
rect 1421 733 1426 737
rect 1419 732 1426 733
rect 1108 726 1121 731
rect 1086 725 1121 726
rect 1141 730 1156 731
rect 1145 726 1156 730
rect 1141 725 1156 726
rect 1158 730 1178 731
rect 1158 726 1174 730
rect 1158 725 1178 726
rect 1185 730 1195 731
rect 1185 726 1187 730
rect 1191 726 1195 730
rect 1185 725 1195 726
rect 1197 730 1216 731
rect 1197 726 1204 730
rect 1208 726 1216 730
rect 1197 725 1216 726
rect 1218 730 1226 731
rect 1218 726 1221 730
rect 1225 726 1226 730
rect 1218 725 1226 726
rect 1239 730 1249 731
rect 1239 726 1241 730
rect 1245 726 1249 730
rect 1239 725 1249 726
rect 1251 730 1270 731
rect 1251 726 1258 730
rect 1262 726 1270 730
rect 1251 725 1270 726
rect 1272 730 1280 731
rect 1272 726 1275 730
rect 1279 726 1280 730
rect 1272 725 1280 726
rect 1295 730 1305 731
rect 1295 726 1297 730
rect 1301 726 1305 730
rect 1295 725 1305 726
rect 1307 730 1326 731
rect 1307 726 1314 730
rect 1318 726 1326 730
rect 1307 725 1326 726
rect 1328 730 1336 731
rect 1328 726 1331 730
rect 1335 726 1336 730
rect 1328 725 1336 726
rect 1349 730 1359 731
rect 1349 726 1351 730
rect 1355 726 1359 730
rect 1349 725 1359 726
rect 1361 730 1380 731
rect 1361 726 1368 730
rect 1372 726 1380 730
rect 1361 725 1380 726
rect 1382 730 1390 731
rect 1382 726 1385 730
rect 1389 726 1390 730
rect 1419 728 1420 732
rect 1424 728 1426 732
rect 1419 727 1426 728
rect 1382 725 1390 726
rect 190 690 198 693
rect 173 685 178 690
rect 171 684 178 685
rect 171 680 172 684
rect 176 680 178 684
rect 171 679 178 680
rect 173 672 178 679
rect 180 672 185 690
rect 187 681 198 690
rect 200 687 205 693
rect 1421 720 1426 727
rect 1428 720 1438 737
rect 1440 741 1445 748
rect 1440 740 1447 741
rect 1440 736 1442 740
rect 1446 736 1447 740
rect 1440 733 1447 736
rect 2071 764 2078 765
rect 2071 760 2072 764
rect 2076 760 2078 764
rect 2071 759 2078 760
rect 2080 785 2092 786
rect 2080 781 2082 785
rect 2086 781 2092 785
rect 2080 778 2092 781
rect 2080 774 2082 778
rect 2086 777 2092 778
rect 2109 777 2114 786
rect 2086 774 2094 777
rect 2080 759 2094 774
rect 2096 764 2104 777
rect 2096 760 2098 764
rect 2102 760 2104 764
rect 2096 759 2104 760
rect 2106 771 2114 777
rect 2106 767 2108 771
rect 2112 767 2114 771
rect 2106 759 2114 767
rect 2116 780 2121 786
rect 2116 779 2123 780
rect 2116 775 2118 779
rect 2122 775 2123 779
rect 2116 774 2123 775
rect 2116 759 2121 774
rect 2157 765 2162 786
rect 2155 764 2162 765
rect 2155 760 2156 764
rect 2160 760 2162 764
rect 2155 759 2162 760
rect 2164 785 2176 786
rect 2164 781 2166 785
rect 2170 781 2176 785
rect 2164 778 2176 781
rect 2164 774 2166 778
rect 2170 777 2176 778
rect 2193 777 2198 786
rect 2170 774 2178 777
rect 2164 759 2178 774
rect 2180 764 2188 777
rect 2180 760 2182 764
rect 2186 760 2188 764
rect 2180 759 2188 760
rect 2190 771 2198 777
rect 2190 767 2192 771
rect 2196 767 2198 771
rect 2190 759 2198 767
rect 2200 780 2205 786
rect 2200 779 2207 780
rect 2200 775 2202 779
rect 2206 775 2207 779
rect 2200 774 2207 775
rect 2200 759 2205 774
rect 2219 764 2224 770
rect 2217 763 2224 764
rect 2217 759 2218 763
rect 2222 759 2224 763
rect 2217 758 2224 759
rect 2226 768 2232 770
rect 2226 763 2234 768
rect 2226 759 2228 763
rect 2232 759 2234 763
rect 2226 758 2234 759
rect 2236 763 2244 768
rect 2236 759 2238 763
rect 2242 759 2244 763
rect 2236 758 2244 759
rect 2246 767 2253 768
rect 2246 763 2248 767
rect 2252 763 2253 767
rect 2246 758 2253 763
rect 1440 729 1442 733
rect 1446 729 1447 733
rect 1440 728 1447 729
rect 1440 720 1445 728
rect 2343 756 2348 762
rect 2341 755 2348 756
rect 2341 751 2342 755
rect 2346 751 2348 755
rect 2341 750 2348 751
rect 2350 760 2356 762
rect 2350 755 2358 760
rect 2350 751 2352 755
rect 2356 751 2358 755
rect 2350 750 2358 751
rect 2360 755 2368 760
rect 2360 751 2362 755
rect 2366 751 2368 755
rect 2360 750 2368 751
rect 2370 759 2377 760
rect 2370 755 2372 759
rect 2376 755 2377 759
rect 2429 757 2434 778
rect 2370 750 2377 755
rect 2427 756 2434 757
rect 2427 752 2428 756
rect 2432 752 2434 756
rect 2427 751 2434 752
rect 2436 777 2448 778
rect 2436 773 2438 777
rect 2442 773 2448 777
rect 2436 770 2448 773
rect 2436 766 2438 770
rect 2442 769 2448 770
rect 2465 769 2470 778
rect 2442 766 2450 769
rect 2436 751 2450 766
rect 2452 756 2460 769
rect 2452 752 2454 756
rect 2458 752 2460 756
rect 2452 751 2460 752
rect 2462 763 2470 769
rect 2462 759 2464 763
rect 2468 759 2470 763
rect 2462 751 2470 759
rect 2472 772 2477 778
rect 2472 771 2479 772
rect 2472 767 2474 771
rect 2478 767 2479 771
rect 2472 766 2479 767
rect 2472 751 2477 766
rect 2513 757 2518 778
rect 2511 756 2518 757
rect 2511 752 2512 756
rect 2516 752 2518 756
rect 2511 751 2518 752
rect 2520 777 2532 778
rect 2520 773 2522 777
rect 2526 773 2532 777
rect 2520 770 2532 773
rect 2520 766 2522 770
rect 2526 769 2532 770
rect 2549 769 2554 778
rect 2526 766 2534 769
rect 2520 751 2534 766
rect 2536 756 2544 769
rect 2536 752 2538 756
rect 2542 752 2544 756
rect 2536 751 2544 752
rect 2546 763 2554 769
rect 2546 759 2548 763
rect 2552 759 2554 763
rect 2546 751 2554 759
rect 2556 772 2561 778
rect 2556 771 2563 772
rect 2556 767 2558 771
rect 2562 767 2563 771
rect 2556 766 2563 767
rect 2556 751 2561 766
rect 2575 756 2580 762
rect 2573 755 2580 756
rect 2573 751 2574 755
rect 2578 751 2580 755
rect 2573 750 2580 751
rect 2582 760 2588 762
rect 2582 755 2590 760
rect 2582 751 2584 755
rect 2588 751 2590 755
rect 2582 750 2590 751
rect 2592 755 2600 760
rect 2592 751 2594 755
rect 2598 751 2600 755
rect 2592 750 2600 751
rect 2602 759 2609 760
rect 2602 755 2604 759
rect 2608 755 2609 759
rect 2703 758 2708 764
rect 2602 750 2609 755
rect 2701 757 2708 758
rect 2701 753 2702 757
rect 2706 753 2708 757
rect 2701 752 2708 753
rect 2710 762 2716 764
rect 2710 757 2718 762
rect 2710 753 2712 757
rect 2716 753 2718 757
rect 2710 752 2718 753
rect 2720 757 2728 762
rect 2720 753 2722 757
rect 2726 753 2728 757
rect 2720 752 2728 753
rect 2730 761 2737 762
rect 2730 757 2732 761
rect 2736 757 2737 761
rect 2789 759 2794 780
rect 2730 752 2737 757
rect 846 695 854 698
rect 519 692 527 695
rect 502 687 507 692
rect 200 686 207 687
rect 200 682 202 686
rect 206 682 207 686
rect 200 681 207 682
rect 500 686 507 687
rect 500 682 501 686
rect 505 682 507 686
rect 500 681 507 682
rect 187 677 196 681
rect 187 673 190 677
rect 194 673 196 677
rect 187 672 196 673
rect 502 674 507 681
rect 509 674 514 692
rect 516 683 527 692
rect 529 689 534 695
rect 829 690 834 695
rect 827 689 834 690
rect 529 688 536 689
rect 529 684 531 688
rect 535 684 536 688
rect 827 685 828 689
rect 832 685 834 689
rect 827 684 834 685
rect 529 683 536 684
rect 516 679 525 683
rect 516 675 519 679
rect 523 675 525 679
rect 829 677 834 684
rect 836 677 841 695
rect 843 686 854 695
rect 856 692 861 698
rect 856 691 863 692
rect 856 687 858 691
rect 862 687 863 691
rect 856 686 863 687
rect 1716 697 1726 698
rect 843 682 852 686
rect 1716 693 1717 697
rect 1721 693 1726 697
rect 1716 691 1726 693
rect 2787 758 2794 759
rect 2787 754 2788 758
rect 2792 754 2794 758
rect 2787 753 2794 754
rect 2796 779 2808 780
rect 2796 775 2798 779
rect 2802 775 2808 779
rect 2796 772 2808 775
rect 2796 768 2798 772
rect 2802 771 2808 772
rect 2825 771 2830 780
rect 2802 768 2810 771
rect 2796 753 2810 768
rect 2812 758 2820 771
rect 2812 754 2814 758
rect 2818 754 2820 758
rect 2812 753 2820 754
rect 2822 765 2830 771
rect 2822 761 2824 765
rect 2828 761 2830 765
rect 2822 753 2830 761
rect 2832 774 2837 780
rect 2832 773 2839 774
rect 2832 769 2834 773
rect 2838 769 2839 773
rect 2832 768 2839 769
rect 2832 753 2837 768
rect 2873 759 2878 780
rect 2871 758 2878 759
rect 2871 754 2872 758
rect 2876 754 2878 758
rect 2871 753 2878 754
rect 2880 779 2892 780
rect 2880 775 2882 779
rect 2886 775 2892 779
rect 2880 772 2892 775
rect 2880 768 2882 772
rect 2886 771 2892 772
rect 2909 771 2914 780
rect 2886 768 2894 771
rect 2880 753 2894 768
rect 2896 758 2904 771
rect 2896 754 2898 758
rect 2902 754 2904 758
rect 2896 753 2904 754
rect 2906 765 2914 771
rect 2906 761 2908 765
rect 2912 761 2914 765
rect 2906 753 2914 761
rect 2916 774 2921 780
rect 2916 773 2923 774
rect 2916 769 2918 773
rect 2922 769 2923 773
rect 2916 768 2923 769
rect 2916 753 2921 768
rect 2935 758 2940 764
rect 2933 757 2940 758
rect 2933 753 2934 757
rect 2938 753 2940 757
rect 2933 752 2940 753
rect 2942 762 2948 764
rect 2942 757 2950 762
rect 2942 753 2944 757
rect 2948 753 2950 757
rect 2942 752 2950 753
rect 2952 757 2960 762
rect 2952 753 2954 757
rect 2958 753 2960 757
rect 2952 752 2960 753
rect 2962 761 2969 762
rect 2962 757 2964 761
rect 2968 757 2969 761
rect 2962 752 2969 757
rect 1716 687 1726 689
rect 843 678 846 682
rect 850 678 852 682
rect 843 677 852 678
rect 516 674 525 675
rect 1716 683 1721 687
rect 1725 683 1726 687
rect 1982 684 1989 685
rect 1716 681 1726 683
rect 1982 680 1983 684
rect 1987 680 1989 684
rect 383 645 389 647
rect 374 640 379 645
rect 372 639 379 640
rect 372 635 373 639
rect 377 635 379 639
rect 372 632 379 635
rect 372 628 373 632
rect 377 628 379 632
rect 372 627 379 628
rect 381 644 389 645
rect 381 640 383 644
rect 387 640 389 644
rect 381 634 389 640
rect 391 646 399 647
rect 391 642 393 646
rect 397 642 399 646
rect 391 639 399 642
rect 391 635 393 639
rect 397 635 399 639
rect 391 634 399 635
rect 401 646 408 647
rect 401 642 403 646
rect 407 642 408 646
rect 476 645 482 647
rect 401 634 408 642
rect 467 640 472 645
rect 465 639 472 640
rect 465 635 466 639
rect 470 635 472 639
rect 381 627 387 634
rect 465 632 472 635
rect 465 628 466 632
rect 470 628 472 632
rect 465 627 472 628
rect 474 644 482 645
rect 474 640 476 644
rect 480 640 482 644
rect 474 634 482 640
rect 484 646 492 647
rect 484 642 486 646
rect 490 642 492 646
rect 484 639 492 642
rect 484 635 486 639
rect 490 635 492 639
rect 484 634 492 635
rect 494 646 501 647
rect 494 642 496 646
rect 500 642 501 646
rect 1650 668 1656 669
rect 1716 677 1726 679
rect 1714 673 1721 677
rect 1725 673 1726 677
rect 1714 671 1726 673
rect 1982 677 1989 680
rect 1982 673 1983 677
rect 1987 673 1989 677
rect 1982 672 1989 673
rect 1650 664 1651 668
rect 1655 667 1656 668
rect 1655 664 1662 667
rect 1650 662 1662 664
rect 1714 667 1726 669
rect 1714 664 1721 667
rect 1720 663 1721 664
rect 1725 663 1726 667
rect 1650 658 1662 660
rect 1650 654 1651 658
rect 1655 654 1662 658
rect 1650 652 1660 654
rect 1720 662 1726 663
rect 1984 657 1989 672
rect 1991 669 1999 685
rect 1991 665 1993 669
rect 1997 665 1999 669
rect 1991 662 1999 665
rect 1991 658 1993 662
rect 1997 658 1999 662
rect 1991 657 1999 658
rect 2001 677 2009 685
rect 2001 673 2003 677
rect 2007 673 2009 677
rect 2001 670 2009 673
rect 2001 666 2003 670
rect 2007 666 2009 670
rect 2001 657 2009 666
rect 2011 669 2022 685
rect 2011 665 2015 669
rect 2019 665 2022 669
rect 2011 662 2022 665
rect 2011 658 2015 662
rect 2019 658 2022 662
rect 2011 657 2022 658
rect 2024 657 2027 685
rect 2029 657 2034 685
rect 2036 682 2041 685
rect 2036 681 2044 682
rect 2036 677 2038 681
rect 2042 677 2044 681
rect 2036 669 2044 677
rect 2046 669 2057 682
rect 2036 657 2041 669
rect 2048 662 2057 669
rect 2048 658 2050 662
rect 2054 658 2057 662
rect 2048 657 2057 658
rect 2059 681 2066 682
rect 2059 677 2061 681
rect 2065 677 2066 681
rect 2059 674 2066 677
rect 2097 674 2105 677
rect 2059 670 2061 674
rect 2065 670 2066 674
rect 2059 669 2066 670
rect 2080 669 2085 674
rect 2059 657 2064 669
rect 2078 668 2085 669
rect 2078 664 2079 668
rect 2083 664 2085 668
rect 2078 663 2085 664
rect 1650 648 1660 650
rect 563 645 569 647
rect 494 634 501 642
rect 554 640 559 645
rect 552 639 559 640
rect 552 635 553 639
rect 557 635 559 639
rect 474 627 480 634
rect 552 632 559 635
rect 552 628 553 632
rect 557 628 559 632
rect 552 627 559 628
rect 561 644 569 645
rect 561 640 563 644
rect 567 640 569 644
rect 561 634 569 640
rect 571 646 579 647
rect 571 642 573 646
rect 577 642 579 646
rect 571 639 579 642
rect 571 635 573 639
rect 577 635 579 639
rect 571 634 579 635
rect 581 646 588 647
rect 581 642 583 646
rect 587 642 588 646
rect 581 634 588 642
rect 561 627 567 634
rect 1650 644 1651 648
rect 1655 644 1660 648
rect 1704 651 1710 652
rect 1704 650 1705 651
rect 1650 642 1660 644
rect 1650 638 1660 640
rect 1650 634 1655 638
rect 1659 634 1660 638
rect 1698 647 1705 650
rect 1709 650 1710 651
rect 1709 647 1725 650
rect 1698 645 1725 647
rect 1698 641 1725 643
rect 1698 638 1713 641
rect 1707 637 1713 638
rect 1717 637 1725 641
rect 1707 635 1725 637
rect 2080 656 2085 663
rect 2087 656 2092 674
rect 2094 665 2105 674
rect 2107 671 2112 677
rect 2107 670 2114 671
rect 2107 666 2109 670
rect 2113 666 2114 670
rect 2453 666 2461 669
rect 2107 665 2114 666
rect 2094 661 2103 665
rect 2436 661 2441 666
rect 2094 657 2097 661
rect 2101 657 2103 661
rect 2434 660 2441 661
rect 2094 656 2103 657
rect 2434 656 2435 660
rect 2439 656 2441 660
rect 2434 655 2441 656
rect 2436 648 2441 655
rect 2443 648 2448 666
rect 2450 657 2461 666
rect 2463 663 2468 669
rect 2813 668 2821 671
rect 2796 663 2801 668
rect 2463 662 2470 663
rect 2463 658 2465 662
rect 2469 658 2470 662
rect 2463 657 2470 658
rect 2794 662 2801 663
rect 2794 658 2795 662
rect 2799 658 2801 662
rect 2794 657 2801 658
rect 2450 653 2459 657
rect 2450 649 2453 653
rect 2457 649 2459 653
rect 2450 648 2459 649
rect 2796 650 2801 657
rect 2803 650 2808 668
rect 2810 659 2821 668
rect 2823 665 2828 671
rect 2823 664 2830 665
rect 2823 660 2825 664
rect 2829 660 2830 664
rect 2823 659 2830 660
rect 2810 655 2819 659
rect 2810 651 2813 655
rect 2817 651 2819 655
rect 2810 650 2819 651
rect 1650 633 1660 634
rect 1145 631 1160 632
rect 1149 627 1160 631
rect 1145 626 1160 627
rect 1162 631 1182 632
rect 1162 627 1178 631
rect 1162 626 1182 627
rect 1189 631 1199 632
rect 1189 627 1191 631
rect 1195 627 1199 631
rect 1189 626 1199 627
rect 1201 631 1220 632
rect 1201 627 1208 631
rect 1212 627 1220 631
rect 1201 626 1220 627
rect 1222 631 1230 632
rect 1222 627 1225 631
rect 1229 627 1230 631
rect 1222 626 1230 627
rect 1243 631 1253 632
rect 1243 627 1245 631
rect 1249 627 1253 631
rect 1243 626 1253 627
rect 1255 631 1274 632
rect 1255 627 1262 631
rect 1266 627 1274 631
rect 1255 626 1274 627
rect 1276 631 1284 632
rect 1276 627 1279 631
rect 1283 627 1284 631
rect 1276 626 1284 627
rect 1299 631 1309 632
rect 1299 627 1301 631
rect 1305 627 1309 631
rect 1299 626 1309 627
rect 1311 631 1330 632
rect 1311 627 1318 631
rect 1322 627 1330 631
rect 1311 626 1330 627
rect 1332 631 1340 632
rect 1332 627 1335 631
rect 1339 627 1340 631
rect 1332 626 1340 627
rect 1353 631 1363 632
rect 1353 627 1355 631
rect 1359 627 1363 631
rect 1353 626 1363 627
rect 1365 631 1384 632
rect 1365 627 1372 631
rect 1376 627 1384 631
rect 1365 626 1384 627
rect 1386 631 1394 632
rect 1386 627 1389 631
rect 1393 627 1394 631
rect 1386 626 1394 627
rect 1707 631 1725 633
rect 1707 627 1720 631
rect 1724 627 1725 631
rect 1707 625 1725 627
rect 1707 621 1725 623
rect 1698 615 1725 621
rect 1698 611 1699 615
rect 1703 611 1706 615
rect 1710 611 1725 615
rect 1698 609 1725 611
rect 1698 605 1725 607
rect 1698 602 1720 605
rect 1719 601 1720 602
rect 1724 601 1725 605
rect 1719 600 1725 601
rect 1555 575 1561 576
rect 1555 574 1556 575
rect 1548 571 1556 574
rect 1560 574 1561 575
rect 1560 571 1566 574
rect 1548 569 1566 571
rect 1548 562 1566 567
rect 1548 557 1566 560
rect 1548 553 1549 557
rect 1553 553 1569 557
rect 1548 551 1569 553
rect 1557 549 1569 551
rect 1557 545 1569 547
rect 1557 541 1558 545
rect 1562 542 1569 545
rect 1562 541 1563 542
rect 1557 540 1563 541
rect 1651 582 1657 583
rect 1651 578 1652 582
rect 1656 581 1657 582
rect 1656 578 1678 581
rect 1651 576 1678 578
rect 1651 572 1678 574
rect 1651 568 1666 572
rect 1670 568 1673 572
rect 1677 568 1678 572
rect 1651 562 1678 568
rect 1704 567 1710 568
rect 1704 566 1705 567
rect 1698 563 1705 566
rect 1709 566 1710 567
rect 1709 563 1725 566
rect 1651 560 1669 562
rect 1698 561 1725 563
rect 1651 556 1669 558
rect 1698 557 1725 559
rect 1651 552 1652 556
rect 1656 552 1669 556
rect 1651 550 1669 552
rect 1698 554 1713 557
rect 1707 553 1713 554
rect 1717 553 1725 557
rect 1707 551 1725 553
rect 1651 546 1669 548
rect 1651 542 1659 546
rect 1663 545 1669 546
rect 1663 542 1678 545
rect 1707 547 1725 549
rect 1707 543 1720 547
rect 1724 543 1725 547
rect 1651 540 1678 542
rect 1707 541 1725 543
rect 1651 536 1678 538
rect 1707 537 1725 539
rect 1651 533 1667 536
rect 1666 532 1667 533
rect 1671 533 1678 536
rect 1671 532 1672 533
rect 1666 531 1672 532
rect 1698 531 1725 537
rect 1698 527 1699 531
rect 1703 527 1706 531
rect 1710 527 1725 531
rect 1698 525 1725 527
rect 1698 521 1725 523
rect 1698 518 1720 521
rect 1719 517 1720 518
rect 1724 517 1725 521
rect 1719 516 1725 517
rect 1813 558 1819 559
rect 1813 557 1814 558
rect 1807 554 1814 557
rect 1818 554 1819 558
rect 1807 552 1819 554
rect 1807 548 1819 550
rect 1807 546 1828 548
rect 1807 542 1823 546
rect 1827 542 1828 546
rect 1810 539 1828 542
rect 1810 532 1828 537
rect 1810 528 1828 530
rect 1810 525 1816 528
rect 1815 524 1816 525
rect 1820 525 1828 528
rect 1820 524 1821 525
rect 1815 523 1821 524
rect 1075 506 1106 507
rect 189 481 195 488
rect 168 473 175 481
rect 168 469 169 473
rect 173 469 175 473
rect 168 468 175 469
rect 177 480 185 481
rect 177 476 179 480
rect 183 476 185 480
rect 177 473 185 476
rect 177 469 179 473
rect 183 469 185 473
rect 177 468 185 469
rect 187 475 195 481
rect 187 471 189 475
rect 193 471 195 475
rect 187 470 195 471
rect 197 487 204 488
rect 197 483 199 487
rect 203 483 204 487
rect 197 480 204 483
rect 276 481 282 488
rect 197 476 199 480
rect 203 476 204 480
rect 197 475 204 476
rect 197 470 202 475
rect 255 473 262 481
rect 187 468 193 470
rect 255 469 256 473
rect 260 469 262 473
rect 255 468 262 469
rect 264 480 272 481
rect 264 476 266 480
rect 270 476 272 480
rect 264 473 272 476
rect 264 469 266 473
rect 270 469 272 473
rect 264 468 272 469
rect 274 475 282 481
rect 274 471 276 475
rect 280 471 282 475
rect 274 470 282 471
rect 284 487 291 488
rect 284 483 286 487
rect 290 483 291 487
rect 284 480 291 483
rect 588 489 595 490
rect 369 481 375 488
rect 284 476 286 480
rect 290 476 291 480
rect 284 475 291 476
rect 284 470 289 475
rect 348 473 355 481
rect 274 468 280 470
rect 348 469 349 473
rect 353 469 355 473
rect 348 468 355 469
rect 357 480 365 481
rect 357 476 359 480
rect 363 476 365 480
rect 357 473 365 476
rect 357 469 359 473
rect 363 469 365 473
rect 357 468 365 469
rect 367 475 375 481
rect 367 471 369 475
rect 373 471 375 475
rect 367 470 375 471
rect 377 487 384 488
rect 377 483 379 487
rect 383 483 384 487
rect 377 480 384 483
rect 377 476 379 480
rect 383 476 384 480
rect 588 485 589 489
rect 593 485 595 489
rect 588 482 595 485
rect 588 478 589 482
rect 593 478 595 482
rect 588 477 595 478
rect 377 475 384 476
rect 377 470 382 475
rect 590 472 595 477
rect 597 483 603 490
rect 681 489 688 490
rect 681 485 682 489
rect 686 485 688 489
rect 597 477 605 483
rect 597 473 599 477
rect 603 473 605 477
rect 597 472 605 473
rect 367 468 373 470
rect 599 470 605 472
rect 607 482 615 483
rect 607 478 609 482
rect 613 478 615 482
rect 607 475 615 478
rect 607 471 609 475
rect 613 471 615 475
rect 607 470 615 471
rect 617 475 624 483
rect 681 482 688 485
rect 681 478 682 482
rect 686 478 688 482
rect 681 477 688 478
rect 617 471 619 475
rect 623 471 624 475
rect 683 472 688 477
rect 690 483 696 490
rect 768 489 775 490
rect 768 485 769 489
rect 773 485 775 489
rect 690 477 698 483
rect 690 473 692 477
rect 696 473 698 477
rect 690 472 698 473
rect 617 470 624 471
rect 692 470 698 472
rect 700 482 708 483
rect 700 478 702 482
rect 706 478 708 482
rect 700 475 708 478
rect 700 471 702 475
rect 706 471 708 475
rect 700 470 708 471
rect 710 475 717 483
rect 768 482 775 485
rect 768 478 769 482
rect 773 478 775 482
rect 768 477 775 478
rect 710 471 712 475
rect 716 471 717 475
rect 770 472 775 477
rect 777 483 783 490
rect 1075 502 1080 506
rect 1084 502 1106 506
rect 1075 501 1106 502
rect 1108 502 1124 507
rect 1130 502 1143 507
rect 1108 501 1143 502
rect 1163 506 1178 507
rect 1167 502 1178 506
rect 1163 501 1178 502
rect 1180 506 1200 507
rect 1180 502 1196 506
rect 1180 501 1200 502
rect 1207 506 1217 507
rect 1207 502 1209 506
rect 1213 502 1217 506
rect 1207 501 1217 502
rect 1219 506 1238 507
rect 1219 502 1226 506
rect 1230 502 1238 506
rect 1219 501 1238 502
rect 1240 506 1248 507
rect 1240 502 1243 506
rect 1247 502 1248 506
rect 1240 501 1248 502
rect 1261 506 1271 507
rect 1261 502 1263 506
rect 1267 502 1271 506
rect 1261 501 1271 502
rect 1273 506 1292 507
rect 1273 502 1280 506
rect 1284 502 1292 506
rect 1273 501 1292 502
rect 1294 506 1302 507
rect 1294 502 1297 506
rect 1301 502 1302 506
rect 1294 501 1302 502
rect 1317 506 1327 507
rect 1317 502 1319 506
rect 1323 502 1327 506
rect 1317 501 1327 502
rect 1329 506 1348 507
rect 1329 502 1336 506
rect 1340 502 1348 506
rect 1329 501 1348 502
rect 1350 506 1358 507
rect 1350 502 1353 506
rect 1357 502 1358 506
rect 1350 501 1358 502
rect 1371 506 1381 507
rect 1371 502 1373 506
rect 1377 502 1381 506
rect 1371 501 1381 502
rect 1383 506 1402 507
rect 1383 502 1390 506
rect 1394 502 1402 506
rect 1383 501 1402 502
rect 1404 506 1412 507
rect 1404 502 1407 506
rect 1411 502 1412 506
rect 1404 501 1412 502
rect 777 477 785 483
rect 777 473 779 477
rect 783 473 785 477
rect 777 472 785 473
rect 710 470 717 471
rect 779 470 785 472
rect 787 482 795 483
rect 787 478 789 482
rect 793 478 795 482
rect 787 475 795 478
rect 787 471 789 475
rect 793 471 795 475
rect 787 470 795 471
rect 797 475 804 483
rect 797 471 799 475
rect 803 471 804 475
rect 797 470 804 471
rect 1651 498 1657 499
rect 1651 494 1652 498
rect 1656 497 1657 498
rect 1656 494 1678 497
rect 1651 492 1678 494
rect 1651 488 1678 490
rect 1651 484 1666 488
rect 1670 484 1673 488
rect 1677 484 1678 488
rect 1651 478 1678 484
rect 1651 476 1669 478
rect 1651 472 1669 474
rect 1651 468 1652 472
rect 1656 468 1669 472
rect 1651 466 1669 468
rect 1716 465 1726 466
rect 1651 462 1669 464
rect 1651 458 1659 462
rect 1663 461 1669 462
rect 1663 458 1678 461
rect 1651 456 1678 458
rect 92 420 97 426
rect 90 419 97 420
rect 90 415 91 419
rect 95 415 97 419
rect 90 414 97 415
rect 99 424 105 426
rect 99 419 107 424
rect 99 415 101 419
rect 105 415 107 419
rect 99 414 107 415
rect 109 419 117 424
rect 109 415 111 419
rect 115 415 117 419
rect 109 414 117 415
rect 119 423 126 424
rect 119 419 121 423
rect 125 419 126 423
rect 178 421 183 442
rect 119 414 126 419
rect 176 420 183 421
rect 176 416 177 420
rect 181 416 183 420
rect 176 415 183 416
rect 185 441 197 442
rect 185 437 187 441
rect 191 437 197 441
rect 185 434 197 437
rect 185 430 187 434
rect 191 433 197 434
rect 214 433 219 442
rect 191 430 199 433
rect 185 415 199 430
rect 201 420 209 433
rect 201 416 203 420
rect 207 416 209 420
rect 201 415 209 416
rect 211 427 219 433
rect 211 423 213 427
rect 217 423 219 427
rect 211 415 219 423
rect 221 436 226 442
rect 221 435 228 436
rect 221 431 223 435
rect 227 431 228 435
rect 221 430 228 431
rect 221 415 226 430
rect 262 421 267 442
rect 260 420 267 421
rect 260 416 261 420
rect 265 416 267 420
rect 260 415 267 416
rect 269 441 281 442
rect 269 437 271 441
rect 275 437 281 441
rect 269 434 281 437
rect 269 430 271 434
rect 275 433 281 434
rect 298 433 303 442
rect 275 430 283 433
rect 269 415 283 430
rect 285 420 293 433
rect 285 416 287 420
rect 291 416 293 420
rect 285 415 293 416
rect 295 427 303 433
rect 295 423 297 427
rect 301 423 303 427
rect 295 415 303 423
rect 305 436 310 442
rect 305 435 312 436
rect 305 431 307 435
rect 311 431 312 435
rect 305 430 312 431
rect 305 415 310 430
rect 324 420 329 426
rect 322 419 329 420
rect 322 415 323 419
rect 327 415 329 419
rect 322 414 329 415
rect 331 424 337 426
rect 331 419 339 424
rect 331 415 333 419
rect 337 415 339 419
rect 331 414 339 415
rect 341 419 349 424
rect 341 415 343 419
rect 347 415 349 419
rect 341 414 349 415
rect 351 423 358 424
rect 351 419 353 423
rect 357 419 358 423
rect 421 422 426 428
rect 351 414 358 419
rect 419 421 426 422
rect 419 417 420 421
rect 424 417 426 421
rect 419 416 426 417
rect 428 426 434 428
rect 428 421 436 426
rect 428 417 430 421
rect 434 417 436 421
rect 428 416 436 417
rect 438 421 446 426
rect 438 417 440 421
rect 444 417 446 421
rect 438 416 446 417
rect 448 425 455 426
rect 448 421 450 425
rect 454 421 455 425
rect 507 423 512 444
rect 448 416 455 421
rect 505 422 512 423
rect 505 418 506 422
rect 510 418 512 422
rect 505 417 512 418
rect 514 443 526 444
rect 514 439 516 443
rect 520 439 526 443
rect 514 436 526 439
rect 514 432 516 436
rect 520 435 526 436
rect 543 435 548 444
rect 520 432 528 435
rect 514 417 528 432
rect 530 422 538 435
rect 530 418 532 422
rect 536 418 538 422
rect 530 417 538 418
rect 540 429 548 435
rect 540 425 542 429
rect 546 425 548 429
rect 540 417 548 425
rect 550 438 555 444
rect 550 437 557 438
rect 550 433 552 437
rect 556 433 557 437
rect 550 432 557 433
rect 550 417 555 432
rect 591 423 596 444
rect 589 422 596 423
rect 589 418 590 422
rect 594 418 596 422
rect 589 417 596 418
rect 598 443 610 444
rect 598 439 600 443
rect 604 439 610 443
rect 598 436 610 439
rect 598 432 600 436
rect 604 435 610 436
rect 627 435 632 444
rect 604 432 612 435
rect 598 417 612 432
rect 614 422 622 435
rect 614 418 616 422
rect 620 418 622 422
rect 614 417 622 418
rect 624 429 632 435
rect 624 425 626 429
rect 630 425 632 429
rect 624 417 632 425
rect 634 438 639 444
rect 634 437 641 438
rect 634 433 636 437
rect 640 433 641 437
rect 634 432 641 433
rect 634 417 639 432
rect 653 422 658 428
rect 651 421 658 422
rect 651 417 652 421
rect 656 417 658 421
rect 651 416 658 417
rect 660 426 666 428
rect 660 421 668 426
rect 660 417 662 421
rect 666 417 668 421
rect 660 416 668 417
rect 670 421 678 426
rect 670 417 672 421
rect 676 417 678 421
rect 670 416 678 417
rect 680 425 687 426
rect 748 425 753 431
rect 680 421 682 425
rect 686 421 687 425
rect 680 416 687 421
rect 746 424 753 425
rect 746 420 747 424
rect 751 420 753 424
rect 746 419 753 420
rect 755 429 761 431
rect 755 424 763 429
rect 755 420 757 424
rect 761 420 763 424
rect 755 419 763 420
rect 765 424 773 429
rect 765 420 767 424
rect 771 420 773 424
rect 765 419 773 420
rect 775 428 782 429
rect 775 424 777 428
rect 781 424 782 428
rect 834 426 839 447
rect 775 419 782 424
rect 832 425 839 426
rect 832 421 833 425
rect 837 421 839 425
rect 832 420 839 421
rect 841 446 853 447
rect 841 442 843 446
rect 847 442 853 446
rect 841 439 853 442
rect 841 435 843 439
rect 847 438 853 439
rect 870 438 875 447
rect 847 435 855 438
rect 841 420 855 435
rect 857 425 865 438
rect 857 421 859 425
rect 863 421 865 425
rect 857 420 865 421
rect 867 432 875 438
rect 867 428 869 432
rect 873 428 875 432
rect 867 420 875 428
rect 877 441 882 447
rect 877 440 884 441
rect 877 436 879 440
rect 883 436 884 440
rect 877 435 884 436
rect 877 420 882 435
rect 918 426 923 447
rect 916 425 923 426
rect 916 421 917 425
rect 921 421 923 425
rect 916 420 923 421
rect 925 446 937 447
rect 925 442 927 446
rect 931 442 937 446
rect 925 439 937 442
rect 925 435 927 439
rect 931 438 937 439
rect 954 438 959 447
rect 931 435 939 438
rect 925 420 939 435
rect 941 425 949 438
rect 941 421 943 425
rect 947 421 949 425
rect 941 420 949 421
rect 951 432 959 438
rect 951 428 953 432
rect 957 428 959 432
rect 951 420 959 428
rect 961 441 966 447
rect 1651 452 1678 454
rect 1651 449 1667 452
rect 1666 448 1667 449
rect 1671 449 1678 452
rect 1716 461 1717 465
rect 1721 461 1726 465
rect 1716 459 1726 461
rect 1716 455 1726 457
rect 1671 448 1672 449
rect 1666 447 1672 448
rect 1716 451 1721 455
rect 1725 451 1726 455
rect 1716 449 1726 451
rect 961 440 968 441
rect 961 436 963 440
rect 967 436 968 440
rect 961 435 968 436
rect 961 420 966 435
rect 980 425 985 431
rect 978 424 985 425
rect 978 420 979 424
rect 983 420 985 424
rect 978 419 985 420
rect 987 429 993 431
rect 987 424 995 429
rect 987 420 989 424
rect 993 420 995 424
rect 987 419 995 420
rect 997 424 1005 429
rect 997 420 999 424
rect 1003 420 1005 424
rect 997 419 1005 420
rect 1007 428 1014 429
rect 1007 424 1009 428
rect 1013 424 1014 428
rect 1650 436 1656 437
rect 1716 445 1726 447
rect 1714 441 1721 445
rect 1725 441 1726 445
rect 1714 439 1726 441
rect 1650 432 1651 436
rect 1655 435 1656 436
rect 1655 432 1662 435
rect 1650 430 1662 432
rect 1714 435 1726 437
rect 1714 432 1721 435
rect 1720 431 1721 432
rect 1725 431 1726 435
rect 1007 419 1014 424
rect 1650 426 1662 428
rect 1650 422 1651 426
rect 1655 422 1662 426
rect 1650 420 1660 422
rect 1720 430 1726 431
rect 1650 416 1660 418
rect 1650 412 1651 416
rect 1655 412 1660 416
rect 1650 410 1660 412
rect 1167 407 1182 408
rect 1171 403 1182 407
rect 1167 402 1182 403
rect 1184 407 1204 408
rect 1184 403 1200 407
rect 1184 402 1204 403
rect 1211 407 1221 408
rect 1211 403 1213 407
rect 1217 403 1221 407
rect 1211 402 1221 403
rect 1223 407 1242 408
rect 1223 403 1230 407
rect 1234 403 1242 407
rect 1223 402 1242 403
rect 1244 407 1252 408
rect 1244 403 1247 407
rect 1251 403 1252 407
rect 1244 402 1252 403
rect 1265 407 1275 408
rect 1265 403 1267 407
rect 1271 403 1275 407
rect 1265 402 1275 403
rect 1277 407 1296 408
rect 1277 403 1284 407
rect 1288 403 1296 407
rect 1277 402 1296 403
rect 1298 407 1306 408
rect 1298 403 1301 407
rect 1305 403 1306 407
rect 1298 402 1306 403
rect 1321 407 1331 408
rect 1321 403 1323 407
rect 1327 403 1331 407
rect 1321 402 1331 403
rect 1333 407 1352 408
rect 1333 403 1340 407
rect 1344 403 1352 407
rect 1333 402 1352 403
rect 1354 407 1362 408
rect 1354 403 1357 407
rect 1361 403 1362 407
rect 1354 402 1362 403
rect 1375 407 1385 408
rect 1375 403 1377 407
rect 1381 403 1385 407
rect 1375 402 1385 403
rect 1387 407 1406 408
rect 1387 403 1394 407
rect 1398 403 1406 407
rect 1387 402 1406 403
rect 1408 407 1416 408
rect 1408 403 1411 407
rect 1415 403 1416 407
rect 1408 402 1416 403
rect 1650 406 1660 408
rect 1650 402 1655 406
rect 1659 402 1660 406
rect 2054 410 2060 417
rect 2033 402 2040 410
rect 1650 401 1660 402
rect 2033 398 2034 402
rect 2038 398 2040 402
rect 2033 397 2040 398
rect 2042 409 2050 410
rect 2042 405 2044 409
rect 2048 405 2050 409
rect 2042 402 2050 405
rect 2042 398 2044 402
rect 2048 398 2050 402
rect 2042 397 2050 398
rect 2052 404 2060 410
rect 2052 400 2054 404
rect 2058 400 2060 404
rect 2052 399 2060 400
rect 2062 416 2069 417
rect 2062 412 2064 416
rect 2068 412 2069 416
rect 2062 409 2069 412
rect 2141 410 2147 417
rect 2062 405 2064 409
rect 2068 405 2069 409
rect 2062 404 2069 405
rect 2062 399 2067 404
rect 2120 402 2127 410
rect 2052 397 2058 399
rect 2120 398 2121 402
rect 2125 398 2127 402
rect 2120 397 2127 398
rect 2129 409 2137 410
rect 2129 405 2131 409
rect 2135 405 2137 409
rect 2129 402 2137 405
rect 2129 398 2131 402
rect 2135 398 2137 402
rect 2129 397 2137 398
rect 2139 404 2147 410
rect 2139 400 2141 404
rect 2145 400 2147 404
rect 2139 399 2147 400
rect 2149 416 2156 417
rect 2149 412 2151 416
rect 2155 412 2156 416
rect 2149 409 2156 412
rect 2453 418 2460 419
rect 2234 410 2240 417
rect 2149 405 2151 409
rect 2155 405 2156 409
rect 2149 404 2156 405
rect 2149 399 2154 404
rect 2213 402 2220 410
rect 2139 397 2145 399
rect 2213 398 2214 402
rect 2218 398 2220 402
rect 2213 397 2220 398
rect 2222 409 2230 410
rect 2222 405 2224 409
rect 2228 405 2230 409
rect 2222 402 2230 405
rect 2222 398 2224 402
rect 2228 398 2230 402
rect 2222 397 2230 398
rect 2232 404 2240 410
rect 2232 400 2234 404
rect 2238 400 2240 404
rect 2232 399 2240 400
rect 2242 416 2249 417
rect 2242 412 2244 416
rect 2248 412 2249 416
rect 2242 409 2249 412
rect 2242 405 2244 409
rect 2248 405 2249 409
rect 2453 414 2454 418
rect 2458 414 2460 418
rect 2453 411 2460 414
rect 2453 407 2454 411
rect 2458 407 2460 411
rect 2453 406 2460 407
rect 2242 404 2249 405
rect 2242 399 2247 404
rect 2455 401 2460 406
rect 2462 412 2468 419
rect 2546 418 2553 419
rect 2546 414 2547 418
rect 2551 414 2553 418
rect 2462 406 2470 412
rect 2462 402 2464 406
rect 2468 402 2470 406
rect 2462 401 2470 402
rect 2232 397 2238 399
rect 2464 399 2470 401
rect 2472 411 2480 412
rect 2472 407 2474 411
rect 2478 407 2480 411
rect 2472 404 2480 407
rect 2472 400 2474 404
rect 2478 400 2480 404
rect 2472 399 2480 400
rect 2482 404 2489 412
rect 2546 411 2553 414
rect 2546 407 2547 411
rect 2551 407 2553 411
rect 2546 406 2553 407
rect 2482 400 2484 404
rect 2488 400 2489 404
rect 2548 401 2553 406
rect 2555 412 2561 419
rect 2633 418 2640 419
rect 2633 414 2634 418
rect 2638 414 2640 418
rect 2555 406 2563 412
rect 2555 402 2557 406
rect 2561 402 2563 406
rect 2555 401 2563 402
rect 2482 399 2489 400
rect 2557 399 2563 401
rect 2565 411 2573 412
rect 2565 407 2567 411
rect 2571 407 2573 411
rect 2565 404 2573 407
rect 2565 400 2567 404
rect 2571 400 2573 404
rect 2565 399 2573 400
rect 2575 404 2582 412
rect 2633 411 2640 414
rect 2633 407 2634 411
rect 2638 407 2640 411
rect 2633 406 2640 407
rect 2575 400 2577 404
rect 2581 400 2582 404
rect 2635 401 2640 406
rect 2642 412 2648 419
rect 2642 406 2650 412
rect 2642 402 2644 406
rect 2648 402 2650 406
rect 2642 401 2650 402
rect 2575 399 2582 400
rect 2644 399 2650 401
rect 2652 411 2660 412
rect 2652 407 2654 411
rect 2658 407 2660 411
rect 2652 404 2660 407
rect 2652 400 2654 404
rect 2658 400 2660 404
rect 2652 399 2660 400
rect 2662 404 2669 412
rect 2662 400 2664 404
rect 2668 400 2669 404
rect 2662 399 2669 400
rect 202 330 210 333
rect 185 325 190 330
rect 183 324 190 325
rect 183 320 184 324
rect 188 320 190 324
rect 183 319 190 320
rect 185 312 190 319
rect 192 312 197 330
rect 199 321 210 330
rect 212 327 217 333
rect 1073 361 1104 362
rect 1073 357 1078 361
rect 1082 357 1104 361
rect 1073 356 1104 357
rect 1106 357 1122 362
rect 1128 357 1141 362
rect 1106 356 1141 357
rect 1161 361 1176 362
rect 1165 357 1176 361
rect 1161 356 1176 357
rect 1178 361 1198 362
rect 1178 357 1194 361
rect 1178 356 1198 357
rect 1205 361 1215 362
rect 1205 357 1207 361
rect 1211 357 1215 361
rect 1205 356 1215 357
rect 1217 361 1236 362
rect 1217 357 1224 361
rect 1228 357 1236 361
rect 1217 356 1236 357
rect 1238 361 1246 362
rect 1238 357 1241 361
rect 1245 357 1246 361
rect 1238 356 1246 357
rect 1259 361 1269 362
rect 1259 357 1261 361
rect 1265 357 1269 361
rect 1259 356 1269 357
rect 1271 361 1290 362
rect 1271 357 1278 361
rect 1282 357 1290 361
rect 1271 356 1290 357
rect 1292 361 1300 362
rect 1292 357 1295 361
rect 1299 357 1300 361
rect 1292 356 1300 357
rect 1315 361 1325 362
rect 1315 357 1317 361
rect 1321 357 1325 361
rect 1315 356 1325 357
rect 1327 361 1346 362
rect 1327 357 1334 361
rect 1338 357 1346 361
rect 1327 356 1346 357
rect 1348 361 1356 362
rect 1348 357 1351 361
rect 1355 357 1356 361
rect 1348 356 1356 357
rect 1369 361 1379 362
rect 1369 357 1371 361
rect 1375 357 1379 361
rect 1369 356 1379 357
rect 1381 361 1400 362
rect 1381 357 1388 361
rect 1392 357 1400 361
rect 1381 356 1400 357
rect 1402 361 1410 362
rect 1402 357 1405 361
rect 1409 357 1410 361
rect 1402 356 1410 357
rect 1957 349 1962 355
rect 858 335 866 338
rect 531 332 539 335
rect 514 327 519 332
rect 212 326 219 327
rect 212 322 214 326
rect 218 322 219 326
rect 212 321 219 322
rect 512 326 519 327
rect 512 322 513 326
rect 517 322 519 326
rect 512 321 519 322
rect 199 317 208 321
rect 199 313 202 317
rect 206 313 208 317
rect 199 312 208 313
rect 514 314 519 321
rect 521 314 526 332
rect 528 323 539 332
rect 541 329 546 335
rect 841 330 846 335
rect 839 329 846 330
rect 541 328 548 329
rect 541 324 543 328
rect 547 324 548 328
rect 839 325 840 329
rect 844 325 846 329
rect 839 324 846 325
rect 541 323 548 324
rect 528 319 537 323
rect 528 315 531 319
rect 535 315 537 319
rect 841 317 846 324
rect 848 317 853 335
rect 855 326 866 335
rect 868 332 873 338
rect 868 331 875 332
rect 868 327 870 331
rect 874 327 875 331
rect 868 326 875 327
rect 855 322 864 326
rect 855 318 858 322
rect 862 318 864 322
rect 1955 348 1962 349
rect 855 317 864 318
rect 528 314 537 315
rect 1955 344 1956 348
rect 1960 344 1962 348
rect 1955 343 1962 344
rect 1964 353 1970 355
rect 1964 348 1972 353
rect 1964 344 1966 348
rect 1970 344 1972 348
rect 1964 343 1972 344
rect 1974 348 1982 353
rect 1974 344 1976 348
rect 1980 344 1982 348
rect 1974 343 1982 344
rect 1984 352 1991 353
rect 1984 348 1986 352
rect 1990 348 1991 352
rect 2043 350 2048 371
rect 1984 343 1991 348
rect 1708 341 1718 342
rect 1708 337 1709 341
rect 1713 337 1718 341
rect 1708 335 1718 337
rect 1708 331 1718 333
rect 1708 327 1713 331
rect 1717 327 1718 331
rect 1708 325 1718 327
rect 1453 307 1458 314
rect 1451 306 1458 307
rect 91 274 96 280
rect 89 273 96 274
rect 89 269 90 273
rect 94 269 96 273
rect 89 268 96 269
rect 98 278 104 280
rect 98 273 106 278
rect 98 269 100 273
rect 104 269 106 273
rect 98 268 106 269
rect 108 273 116 278
rect 108 269 110 273
rect 114 269 116 273
rect 108 268 116 269
rect 118 277 125 278
rect 118 273 120 277
rect 124 273 125 277
rect 177 275 182 296
rect 118 268 125 273
rect 175 274 182 275
rect 175 270 176 274
rect 180 270 182 274
rect 175 269 182 270
rect 184 295 196 296
rect 184 291 186 295
rect 190 291 196 295
rect 184 288 196 291
rect 184 284 186 288
rect 190 287 196 288
rect 213 287 218 296
rect 190 284 198 287
rect 184 269 198 284
rect 200 274 208 287
rect 200 270 202 274
rect 206 270 208 274
rect 200 269 208 270
rect 210 281 218 287
rect 210 277 212 281
rect 216 277 218 281
rect 210 269 218 277
rect 220 290 225 296
rect 220 289 227 290
rect 220 285 222 289
rect 226 285 227 289
rect 220 284 227 285
rect 220 269 225 284
rect 261 275 266 296
rect 259 274 266 275
rect 259 270 260 274
rect 264 270 266 274
rect 259 269 266 270
rect 268 295 280 296
rect 268 291 270 295
rect 274 291 280 295
rect 268 288 280 291
rect 268 284 270 288
rect 274 287 280 288
rect 297 287 302 296
rect 274 284 282 287
rect 268 269 282 284
rect 284 274 292 287
rect 284 270 286 274
rect 290 270 292 274
rect 284 269 292 270
rect 294 281 302 287
rect 294 277 296 281
rect 300 277 302 281
rect 294 269 302 277
rect 304 290 309 296
rect 304 289 311 290
rect 304 285 306 289
rect 310 285 311 289
rect 304 284 311 285
rect 304 269 309 284
rect 323 274 328 280
rect 321 273 328 274
rect 321 269 322 273
rect 326 269 328 273
rect 321 268 328 269
rect 330 278 336 280
rect 330 273 338 278
rect 330 269 332 273
rect 336 269 338 273
rect 330 268 338 269
rect 340 273 348 278
rect 340 269 342 273
rect 346 269 348 273
rect 340 268 348 269
rect 350 277 357 278
rect 350 273 352 277
rect 356 273 357 277
rect 420 276 425 282
rect 350 268 357 273
rect 418 275 425 276
rect 418 271 419 275
rect 423 271 425 275
rect 418 270 425 271
rect 427 280 433 282
rect 427 275 435 280
rect 427 271 429 275
rect 433 271 435 275
rect 427 270 435 271
rect 437 275 445 280
rect 437 271 439 275
rect 443 271 445 275
rect 437 270 445 271
rect 447 279 454 280
rect 447 275 449 279
rect 453 275 454 279
rect 506 277 511 298
rect 447 270 454 275
rect 504 276 511 277
rect 504 272 505 276
rect 509 272 511 276
rect 504 271 511 272
rect 513 297 525 298
rect 513 293 515 297
rect 519 293 525 297
rect 513 290 525 293
rect 513 286 515 290
rect 519 289 525 290
rect 542 289 547 298
rect 519 286 527 289
rect 513 271 527 286
rect 529 276 537 289
rect 529 272 531 276
rect 535 272 537 276
rect 529 271 537 272
rect 539 283 547 289
rect 539 279 541 283
rect 545 279 547 283
rect 539 271 547 279
rect 549 292 554 298
rect 549 291 556 292
rect 549 287 551 291
rect 555 287 556 291
rect 549 286 556 287
rect 549 271 554 286
rect 590 277 595 298
rect 588 276 595 277
rect 588 272 589 276
rect 593 272 595 276
rect 588 271 595 272
rect 597 297 609 298
rect 597 293 599 297
rect 603 293 609 297
rect 597 290 609 293
rect 597 286 599 290
rect 603 289 609 290
rect 626 289 631 298
rect 603 286 611 289
rect 597 271 611 286
rect 613 276 621 289
rect 613 272 615 276
rect 619 272 621 276
rect 613 271 621 272
rect 623 283 631 289
rect 623 279 625 283
rect 629 279 631 283
rect 623 271 631 279
rect 633 292 638 298
rect 633 291 640 292
rect 633 287 635 291
rect 639 287 640 291
rect 633 286 640 287
rect 633 271 638 286
rect 652 276 657 282
rect 650 275 657 276
rect 650 271 651 275
rect 655 271 657 275
rect 650 270 657 271
rect 659 280 665 282
rect 659 275 667 280
rect 659 271 661 275
rect 665 271 667 275
rect 659 270 667 271
rect 669 275 677 280
rect 669 271 671 275
rect 675 271 677 275
rect 669 270 677 271
rect 679 279 686 280
rect 747 279 752 285
rect 679 275 681 279
rect 685 275 686 279
rect 679 270 686 275
rect 745 278 752 279
rect 745 274 746 278
rect 750 274 752 278
rect 745 273 752 274
rect 754 283 760 285
rect 754 278 762 283
rect 754 274 756 278
rect 760 274 762 278
rect 754 273 762 274
rect 764 278 772 283
rect 764 274 766 278
rect 770 274 772 278
rect 764 273 772 274
rect 774 282 781 283
rect 774 278 776 282
rect 780 278 781 282
rect 833 280 838 301
rect 774 273 781 278
rect 831 279 838 280
rect 831 275 832 279
rect 836 275 838 279
rect 831 274 838 275
rect 840 300 852 301
rect 840 296 842 300
rect 846 296 852 300
rect 840 293 852 296
rect 840 289 842 293
rect 846 292 852 293
rect 869 292 874 301
rect 846 289 854 292
rect 840 274 854 289
rect 856 279 864 292
rect 856 275 858 279
rect 862 275 864 279
rect 856 274 864 275
rect 866 286 874 292
rect 866 282 868 286
rect 872 282 874 286
rect 866 274 874 282
rect 876 295 881 301
rect 876 294 883 295
rect 876 290 878 294
rect 882 290 883 294
rect 876 289 883 290
rect 876 274 881 289
rect 917 280 922 301
rect 915 279 922 280
rect 915 275 916 279
rect 920 275 922 279
rect 915 274 922 275
rect 924 300 936 301
rect 924 296 926 300
rect 930 296 936 300
rect 924 293 936 296
rect 924 289 926 293
rect 930 292 936 293
rect 953 292 958 301
rect 930 289 938 292
rect 924 274 938 289
rect 940 279 948 292
rect 940 275 942 279
rect 946 275 948 279
rect 940 274 948 275
rect 950 286 958 292
rect 950 282 952 286
rect 956 282 958 286
rect 950 274 958 282
rect 960 295 965 301
rect 1451 302 1452 306
rect 1456 302 1458 306
rect 1451 301 1458 302
rect 960 294 967 295
rect 960 290 962 294
rect 966 290 967 294
rect 960 289 967 290
rect 960 274 965 289
rect 979 279 984 285
rect 977 278 984 279
rect 977 274 978 278
rect 982 274 984 278
rect 977 273 984 274
rect 986 283 992 285
rect 986 278 994 283
rect 986 274 988 278
rect 992 274 994 278
rect 986 273 994 274
rect 996 278 1004 283
rect 996 274 998 278
rect 1002 274 1004 278
rect 996 273 1004 274
rect 1006 282 1013 283
rect 1006 278 1008 282
rect 1012 278 1013 282
rect 1453 297 1458 301
rect 1460 297 1470 314
rect 1462 288 1470 297
rect 1462 284 1463 288
rect 1467 286 1470 288
rect 1472 306 1477 314
rect 1708 321 1718 323
rect 1706 317 1713 321
rect 1717 317 1718 321
rect 1706 315 1718 317
rect 2041 349 2048 350
rect 2041 345 2042 349
rect 2046 345 2048 349
rect 2041 344 2048 345
rect 2050 370 2062 371
rect 2050 366 2052 370
rect 2056 366 2062 370
rect 2050 363 2062 366
rect 2050 359 2052 363
rect 2056 362 2062 363
rect 2079 362 2084 371
rect 2056 359 2064 362
rect 2050 344 2064 359
rect 2066 349 2074 362
rect 2066 345 2068 349
rect 2072 345 2074 349
rect 2066 344 2074 345
rect 2076 356 2084 362
rect 2076 352 2078 356
rect 2082 352 2084 356
rect 2076 344 2084 352
rect 2086 365 2091 371
rect 2086 364 2093 365
rect 2086 360 2088 364
rect 2092 360 2093 364
rect 2086 359 2093 360
rect 2086 344 2091 359
rect 2127 350 2132 371
rect 2125 349 2132 350
rect 2125 345 2126 349
rect 2130 345 2132 349
rect 2125 344 2132 345
rect 2134 370 2146 371
rect 2134 366 2136 370
rect 2140 366 2146 370
rect 2134 363 2146 366
rect 2134 359 2136 363
rect 2140 362 2146 363
rect 2163 362 2168 371
rect 2140 359 2148 362
rect 2134 344 2148 359
rect 2150 349 2158 362
rect 2150 345 2152 349
rect 2156 345 2158 349
rect 2150 344 2158 345
rect 2160 356 2168 362
rect 2160 352 2162 356
rect 2166 352 2168 356
rect 2160 344 2168 352
rect 2170 365 2175 371
rect 2170 364 2177 365
rect 2170 360 2172 364
rect 2176 360 2177 364
rect 2170 359 2177 360
rect 2170 344 2175 359
rect 2189 349 2194 355
rect 2187 348 2194 349
rect 2187 344 2188 348
rect 2192 344 2194 348
rect 2187 343 2194 344
rect 2196 353 2202 355
rect 2196 348 2204 353
rect 2196 344 2198 348
rect 2202 344 2204 348
rect 2196 343 2204 344
rect 2206 348 2214 353
rect 2206 344 2208 348
rect 2212 344 2214 348
rect 2206 343 2214 344
rect 2216 352 2223 353
rect 2216 348 2218 352
rect 2222 348 2223 352
rect 2286 351 2291 357
rect 2216 343 2223 348
rect 2284 350 2291 351
rect 2284 346 2285 350
rect 2289 346 2291 350
rect 2284 345 2291 346
rect 2293 355 2299 357
rect 2293 350 2301 355
rect 2293 346 2295 350
rect 2299 346 2301 350
rect 2293 345 2301 346
rect 2303 350 2311 355
rect 2303 346 2305 350
rect 2309 346 2311 350
rect 2303 345 2311 346
rect 2313 354 2320 355
rect 2313 350 2315 354
rect 2319 350 2320 354
rect 2372 352 2377 373
rect 2313 345 2320 350
rect 1706 311 1718 313
rect 1706 308 1713 311
rect 1712 307 1713 308
rect 1717 307 1718 311
rect 1712 306 1718 307
rect 2370 351 2377 352
rect 2370 347 2371 351
rect 2375 347 2377 351
rect 2370 346 2377 347
rect 2379 372 2391 373
rect 2379 368 2381 372
rect 2385 368 2391 372
rect 2379 365 2391 368
rect 2379 361 2381 365
rect 2385 364 2391 365
rect 2408 364 2413 373
rect 2385 361 2393 364
rect 2379 346 2393 361
rect 2395 351 2403 364
rect 2395 347 2397 351
rect 2401 347 2403 351
rect 2395 346 2403 347
rect 2405 358 2413 364
rect 2405 354 2407 358
rect 2411 354 2413 358
rect 2405 346 2413 354
rect 2415 367 2420 373
rect 2415 366 2422 367
rect 2415 362 2417 366
rect 2421 362 2422 366
rect 2415 361 2422 362
rect 2415 346 2420 361
rect 2456 352 2461 373
rect 2454 351 2461 352
rect 2454 347 2455 351
rect 2459 347 2461 351
rect 2454 346 2461 347
rect 2463 372 2475 373
rect 2463 368 2465 372
rect 2469 368 2475 372
rect 2463 365 2475 368
rect 2463 361 2465 365
rect 2469 364 2475 365
rect 2492 364 2497 373
rect 2469 361 2477 364
rect 2463 346 2477 361
rect 2479 351 2487 364
rect 2479 347 2481 351
rect 2485 347 2487 351
rect 2479 346 2487 347
rect 2489 358 2497 364
rect 2489 354 2491 358
rect 2495 354 2497 358
rect 2489 346 2497 354
rect 2499 367 2504 373
rect 2499 366 2506 367
rect 2499 362 2501 366
rect 2505 362 2506 366
rect 2499 361 2506 362
rect 2499 346 2504 361
rect 2518 351 2523 357
rect 2516 350 2523 351
rect 2516 346 2517 350
rect 2521 346 2523 350
rect 2516 345 2523 346
rect 2525 355 2531 357
rect 2525 350 2533 355
rect 2525 346 2527 350
rect 2531 346 2533 350
rect 2525 345 2533 346
rect 2535 350 2543 355
rect 2535 346 2537 350
rect 2541 346 2543 350
rect 2535 345 2543 346
rect 2545 354 2552 355
rect 2613 354 2618 360
rect 2545 350 2547 354
rect 2551 350 2552 354
rect 2545 345 2552 350
rect 2611 353 2618 354
rect 2611 349 2612 353
rect 2616 349 2618 353
rect 2611 348 2618 349
rect 2620 358 2626 360
rect 2620 353 2628 358
rect 2620 349 2622 353
rect 2626 349 2628 353
rect 2620 348 2628 349
rect 2630 353 2638 358
rect 2630 349 2632 353
rect 2636 349 2638 353
rect 2630 348 2638 349
rect 2640 357 2647 358
rect 2640 353 2642 357
rect 2646 353 2647 357
rect 2699 355 2704 376
rect 2640 348 2647 353
rect 2697 354 2704 355
rect 2697 350 2698 354
rect 2702 350 2704 354
rect 2697 349 2704 350
rect 2706 375 2718 376
rect 2706 371 2708 375
rect 2712 371 2718 375
rect 2706 368 2718 371
rect 2706 364 2708 368
rect 2712 367 2718 368
rect 2735 367 2740 376
rect 2712 364 2720 367
rect 2706 349 2720 364
rect 2722 354 2730 367
rect 2722 350 2724 354
rect 2728 350 2730 354
rect 2722 349 2730 350
rect 2732 361 2740 367
rect 2732 357 2734 361
rect 2738 357 2740 361
rect 2732 349 2740 357
rect 2742 370 2747 376
rect 2742 369 2749 370
rect 2742 365 2744 369
rect 2748 365 2749 369
rect 2742 364 2749 365
rect 2742 349 2747 364
rect 2783 355 2788 376
rect 2781 354 2788 355
rect 2781 350 2782 354
rect 2786 350 2788 354
rect 2781 349 2788 350
rect 2790 375 2802 376
rect 2790 371 2792 375
rect 2796 371 2802 375
rect 2790 368 2802 371
rect 2790 364 2792 368
rect 2796 367 2802 368
rect 2819 367 2824 376
rect 2796 364 2804 367
rect 2790 349 2804 364
rect 2806 354 2814 367
rect 2806 350 2808 354
rect 2812 350 2814 354
rect 2806 349 2814 350
rect 2816 361 2824 367
rect 2816 357 2818 361
rect 2822 357 2824 361
rect 2816 349 2824 357
rect 2826 370 2831 376
rect 2826 369 2833 370
rect 2826 365 2828 369
rect 2832 365 2833 369
rect 2826 364 2833 365
rect 2826 349 2831 364
rect 2845 354 2850 360
rect 2843 353 2850 354
rect 2843 349 2844 353
rect 2848 349 2850 353
rect 2843 348 2850 349
rect 2852 358 2858 360
rect 2852 353 2860 358
rect 2852 349 2854 353
rect 2858 349 2860 353
rect 2852 348 2860 349
rect 2862 353 2870 358
rect 2862 349 2864 353
rect 2868 349 2870 353
rect 2862 348 2870 349
rect 2872 357 2879 358
rect 2872 353 2874 357
rect 2878 353 2879 357
rect 2872 348 2879 353
rect 1472 305 1479 306
rect 1472 301 1474 305
rect 1478 301 1479 305
rect 1472 298 1479 301
rect 1472 294 1474 298
rect 1478 294 1479 298
rect 1696 295 1702 296
rect 1696 294 1697 295
rect 1472 293 1479 294
rect 1472 286 1477 293
rect 1690 291 1697 294
rect 1701 294 1702 295
rect 1701 291 1717 294
rect 1690 289 1717 291
rect 1467 284 1468 286
rect 1462 283 1468 284
rect 1690 285 1717 287
rect 1690 282 1705 285
rect 1699 281 1705 282
rect 1709 281 1717 285
rect 1699 279 1717 281
rect 1006 273 1013 278
rect 1699 275 1717 277
rect 1699 271 1712 275
rect 1716 271 1717 275
rect 1699 269 1717 271
rect 1699 265 1717 267
rect 1165 262 1180 263
rect 1169 258 1180 262
rect 1165 257 1180 258
rect 1182 262 1202 263
rect 1182 258 1198 262
rect 1182 257 1202 258
rect 1209 262 1219 263
rect 1209 258 1211 262
rect 1215 258 1219 262
rect 1209 257 1219 258
rect 1221 262 1240 263
rect 1221 258 1228 262
rect 1232 258 1240 262
rect 1221 257 1240 258
rect 1242 262 1250 263
rect 1242 258 1245 262
rect 1249 258 1250 262
rect 1242 257 1250 258
rect 1263 262 1273 263
rect 1263 258 1265 262
rect 1269 258 1273 262
rect 1263 257 1273 258
rect 1275 262 1294 263
rect 1275 258 1282 262
rect 1286 258 1294 262
rect 1275 257 1294 258
rect 1296 262 1304 263
rect 1296 258 1299 262
rect 1303 258 1304 262
rect 1296 257 1304 258
rect 1319 262 1329 263
rect 1319 258 1321 262
rect 1325 258 1329 262
rect 1319 257 1329 258
rect 1331 262 1350 263
rect 1331 258 1338 262
rect 1342 258 1350 262
rect 1331 257 1350 258
rect 1352 262 1360 263
rect 1352 258 1355 262
rect 1359 258 1360 262
rect 1352 257 1360 258
rect 1373 262 1383 263
rect 1373 258 1375 262
rect 1379 258 1383 262
rect 1373 257 1383 258
rect 1385 262 1404 263
rect 1385 258 1392 262
rect 1396 258 1404 262
rect 1385 257 1404 258
rect 1406 262 1414 263
rect 1406 258 1409 262
rect 1413 258 1414 262
rect 1406 257 1414 258
rect 1690 259 1717 265
rect 1464 255 1470 256
rect 1464 251 1465 255
rect 1469 253 1470 255
rect 1690 255 1691 259
rect 1695 255 1698 259
rect 1702 255 1717 259
rect 1690 253 1717 255
rect 1469 251 1472 253
rect 1464 242 1472 251
rect 1455 238 1460 242
rect 1453 237 1460 238
rect 1453 233 1454 237
rect 1458 233 1460 237
rect 1453 232 1460 233
rect 1074 219 1105 220
rect 201 184 209 187
rect 184 179 189 184
rect 182 178 189 179
rect 182 174 183 178
rect 187 174 189 178
rect 182 173 189 174
rect 184 166 189 173
rect 191 166 196 184
rect 198 175 209 184
rect 211 181 216 187
rect 1074 215 1079 219
rect 1083 215 1105 219
rect 1074 214 1105 215
rect 1107 215 1123 220
rect 1455 225 1460 232
rect 1462 225 1472 242
rect 1474 246 1479 253
rect 1690 249 1717 251
rect 1690 246 1712 249
rect 1474 245 1481 246
rect 1474 241 1476 245
rect 1480 241 1481 245
rect 1711 245 1712 246
rect 1716 245 1717 249
rect 1711 244 1717 245
rect 2067 259 2075 262
rect 2050 254 2055 259
rect 2048 253 2055 254
rect 2048 249 2049 253
rect 2053 249 2055 253
rect 2048 248 2055 249
rect 1474 238 1481 241
rect 1474 234 1476 238
rect 1480 234 1481 238
rect 2050 241 2055 248
rect 2057 241 2062 259
rect 2064 250 2075 259
rect 2077 256 2082 262
rect 2723 264 2731 267
rect 2396 261 2404 264
rect 2379 256 2384 261
rect 2077 255 2084 256
rect 2077 251 2079 255
rect 2083 251 2084 255
rect 2077 250 2084 251
rect 2377 255 2384 256
rect 2377 251 2378 255
rect 2382 251 2384 255
rect 2377 250 2384 251
rect 2064 246 2073 250
rect 2064 242 2067 246
rect 2071 242 2073 246
rect 2064 241 2073 242
rect 2379 243 2384 250
rect 2386 243 2391 261
rect 2393 252 2404 261
rect 2406 258 2411 264
rect 2706 259 2711 264
rect 2704 258 2711 259
rect 2406 257 2413 258
rect 2406 253 2408 257
rect 2412 253 2413 257
rect 2704 254 2705 258
rect 2709 254 2711 258
rect 2704 253 2711 254
rect 2406 252 2413 253
rect 2393 248 2402 252
rect 2393 244 2396 248
rect 2400 244 2402 248
rect 2706 246 2711 253
rect 2713 246 2718 264
rect 2720 255 2731 264
rect 2733 261 2738 267
rect 2733 260 2740 261
rect 2733 256 2735 260
rect 2739 256 2740 260
rect 2733 255 2740 256
rect 2720 251 2729 255
rect 2720 247 2723 251
rect 2727 247 2729 251
rect 2720 246 2729 247
rect 2393 243 2402 244
rect 1474 233 1481 234
rect 1474 225 1479 233
rect 1129 215 1142 220
rect 1107 214 1142 215
rect 1162 219 1177 220
rect 1166 215 1177 219
rect 1162 214 1177 215
rect 1179 219 1199 220
rect 1179 215 1195 219
rect 1179 214 1199 215
rect 1206 219 1216 220
rect 1206 215 1208 219
rect 1212 215 1216 219
rect 1206 214 1216 215
rect 1218 219 1237 220
rect 1218 215 1225 219
rect 1229 215 1237 219
rect 1218 214 1237 215
rect 1239 219 1247 220
rect 1239 215 1242 219
rect 1246 215 1247 219
rect 1239 214 1247 215
rect 1260 219 1270 220
rect 1260 215 1262 219
rect 1266 215 1270 219
rect 1260 214 1270 215
rect 1272 219 1291 220
rect 1272 215 1279 219
rect 1283 215 1291 219
rect 1272 214 1291 215
rect 1293 219 1301 220
rect 1293 215 1296 219
rect 1300 215 1301 219
rect 1293 214 1301 215
rect 1316 219 1326 220
rect 1316 215 1318 219
rect 1322 215 1326 219
rect 1316 214 1326 215
rect 1328 219 1347 220
rect 1328 215 1335 219
rect 1339 215 1347 219
rect 1328 214 1347 215
rect 1349 219 1357 220
rect 1349 215 1352 219
rect 1356 215 1357 219
rect 1349 214 1357 215
rect 1370 219 1380 220
rect 1370 215 1372 219
rect 1376 215 1380 219
rect 1370 214 1380 215
rect 1382 219 1401 220
rect 1382 215 1389 219
rect 1393 215 1401 219
rect 1382 214 1401 215
rect 1403 219 1411 220
rect 1403 215 1406 219
rect 1410 215 1411 219
rect 1403 214 1411 215
rect 857 189 865 192
rect 530 186 538 189
rect 513 181 518 186
rect 211 180 218 181
rect 211 176 213 180
rect 217 176 218 180
rect 211 175 218 176
rect 511 180 518 181
rect 511 176 512 180
rect 516 176 518 180
rect 511 175 518 176
rect 198 171 207 175
rect 198 167 201 171
rect 205 167 207 171
rect 198 166 207 167
rect 513 168 518 175
rect 520 168 525 186
rect 527 177 538 186
rect 540 183 545 189
rect 840 184 845 189
rect 838 183 845 184
rect 540 182 547 183
rect 540 178 542 182
rect 546 178 547 182
rect 838 179 839 183
rect 843 179 845 183
rect 838 178 845 179
rect 540 177 547 178
rect 527 173 536 177
rect 527 169 530 173
rect 534 169 536 173
rect 840 171 845 178
rect 847 171 852 189
rect 854 180 865 189
rect 867 186 872 192
rect 867 185 874 186
rect 867 181 869 185
rect 873 181 874 185
rect 867 180 874 181
rect 854 176 863 180
rect 1696 211 1702 212
rect 1696 210 1697 211
rect 1690 207 1697 210
rect 1701 210 1702 211
rect 1701 207 1717 210
rect 1690 205 1717 207
rect 1690 201 1717 203
rect 854 172 857 176
rect 861 172 863 176
rect 1690 198 1705 201
rect 1699 197 1705 198
rect 1709 197 1717 201
rect 1956 203 1961 209
rect 1699 195 1717 197
rect 1699 191 1717 193
rect 1699 187 1712 191
rect 1716 187 1717 191
rect 1699 185 1717 187
rect 1699 181 1717 183
rect 1690 175 1717 181
rect 854 171 863 172
rect 527 168 536 169
rect 1690 171 1691 175
rect 1695 171 1698 175
rect 1702 171 1717 175
rect 1690 169 1717 171
rect 394 139 400 141
rect 385 134 390 139
rect 383 133 390 134
rect 383 129 384 133
rect 388 129 390 133
rect 383 126 390 129
rect 383 122 384 126
rect 388 122 390 126
rect 383 121 390 122
rect 392 138 400 139
rect 392 134 394 138
rect 398 134 400 138
rect 392 128 400 134
rect 402 140 410 141
rect 402 136 404 140
rect 408 136 410 140
rect 402 133 410 136
rect 402 129 404 133
rect 408 129 410 133
rect 402 128 410 129
rect 412 140 419 141
rect 412 136 414 140
rect 418 136 419 140
rect 487 139 493 141
rect 412 128 419 136
rect 478 134 483 139
rect 476 133 483 134
rect 476 129 477 133
rect 481 129 483 133
rect 392 121 398 128
rect 476 126 483 129
rect 476 122 477 126
rect 481 122 483 126
rect 476 121 483 122
rect 485 138 493 139
rect 485 134 487 138
rect 491 134 493 138
rect 485 128 493 134
rect 495 140 503 141
rect 495 136 497 140
rect 501 136 503 140
rect 495 133 503 136
rect 495 129 497 133
rect 501 129 503 133
rect 495 128 503 129
rect 505 140 512 141
rect 505 136 507 140
rect 511 136 512 140
rect 574 139 580 141
rect 505 128 512 136
rect 565 134 570 139
rect 563 133 570 134
rect 563 129 564 133
rect 568 129 570 133
rect 485 121 491 128
rect 563 126 570 129
rect 563 122 564 126
rect 568 122 570 126
rect 563 121 570 122
rect 572 138 580 139
rect 572 134 574 138
rect 578 134 580 138
rect 572 128 580 134
rect 582 140 590 141
rect 582 136 584 140
rect 588 136 590 140
rect 582 133 590 136
rect 582 129 584 133
rect 588 129 590 133
rect 582 128 590 129
rect 592 140 599 141
rect 592 136 594 140
rect 598 136 599 140
rect 1690 165 1717 167
rect 1690 162 1712 165
rect 1711 161 1712 162
rect 1716 161 1717 165
rect 1711 160 1717 161
rect 1805 202 1811 203
rect 1954 202 1961 203
rect 1805 201 1806 202
rect 1799 198 1806 201
rect 1810 198 1811 202
rect 1799 196 1811 198
rect 1954 198 1955 202
rect 1959 198 1961 202
rect 1954 197 1961 198
rect 1963 207 1969 209
rect 1963 202 1971 207
rect 1963 198 1965 202
rect 1969 198 1971 202
rect 1963 197 1971 198
rect 1973 202 1981 207
rect 1973 198 1975 202
rect 1979 198 1981 202
rect 1973 197 1981 198
rect 1983 206 1990 207
rect 1983 202 1985 206
rect 1989 202 1990 206
rect 2042 204 2047 225
rect 1983 197 1990 202
rect 1799 192 1811 194
rect 1799 190 1820 192
rect 1799 186 1815 190
rect 1819 186 1820 190
rect 1802 183 1820 186
rect 1802 176 1820 181
rect 2040 203 2047 204
rect 2040 199 2041 203
rect 2045 199 2047 203
rect 2040 198 2047 199
rect 2049 224 2061 225
rect 2049 220 2051 224
rect 2055 220 2061 224
rect 2049 217 2061 220
rect 2049 213 2051 217
rect 2055 216 2061 217
rect 2078 216 2083 225
rect 2055 213 2063 216
rect 2049 198 2063 213
rect 2065 203 2073 216
rect 2065 199 2067 203
rect 2071 199 2073 203
rect 2065 198 2073 199
rect 2075 210 2083 216
rect 2075 206 2077 210
rect 2081 206 2083 210
rect 2075 198 2083 206
rect 2085 219 2090 225
rect 2085 218 2092 219
rect 2085 214 2087 218
rect 2091 214 2092 218
rect 2085 213 2092 214
rect 2085 198 2090 213
rect 2126 204 2131 225
rect 2124 203 2131 204
rect 2124 199 2125 203
rect 2129 199 2131 203
rect 2124 198 2131 199
rect 2133 224 2145 225
rect 2133 220 2135 224
rect 2139 220 2145 224
rect 2133 217 2145 220
rect 2133 213 2135 217
rect 2139 216 2145 217
rect 2162 216 2167 225
rect 2139 213 2147 216
rect 2133 198 2147 213
rect 2149 203 2157 216
rect 2149 199 2151 203
rect 2155 199 2157 203
rect 2149 198 2157 199
rect 2159 210 2167 216
rect 2159 206 2161 210
rect 2165 206 2167 210
rect 2159 198 2167 206
rect 2169 219 2174 225
rect 2169 218 2176 219
rect 2169 214 2171 218
rect 2175 214 2176 218
rect 2169 213 2176 214
rect 2169 198 2174 213
rect 2188 203 2193 209
rect 2186 202 2193 203
rect 2186 198 2187 202
rect 2191 198 2193 202
rect 2186 197 2193 198
rect 2195 207 2201 209
rect 2195 202 2203 207
rect 2195 198 2197 202
rect 2201 198 2203 202
rect 2195 197 2203 198
rect 2205 202 2213 207
rect 2205 198 2207 202
rect 2211 198 2213 202
rect 2205 197 2213 198
rect 2215 206 2222 207
rect 2215 202 2217 206
rect 2221 202 2222 206
rect 2285 205 2290 211
rect 2215 197 2222 202
rect 2283 204 2290 205
rect 2283 200 2284 204
rect 2288 200 2290 204
rect 2283 199 2290 200
rect 2292 209 2298 211
rect 2292 204 2300 209
rect 2292 200 2294 204
rect 2298 200 2300 204
rect 2292 199 2300 200
rect 2302 204 2310 209
rect 2302 200 2304 204
rect 2308 200 2310 204
rect 2302 199 2310 200
rect 2312 208 2319 209
rect 2312 204 2314 208
rect 2318 204 2319 208
rect 2371 206 2376 227
rect 2312 199 2319 204
rect 1802 172 1820 174
rect 1802 169 1808 172
rect 1807 168 1808 169
rect 1812 169 1820 172
rect 1812 168 1813 169
rect 1807 167 1813 168
rect 2369 205 2376 206
rect 2369 201 2370 205
rect 2374 201 2376 205
rect 2369 200 2376 201
rect 2378 226 2390 227
rect 2378 222 2380 226
rect 2384 222 2390 226
rect 2378 219 2390 222
rect 2378 215 2380 219
rect 2384 218 2390 219
rect 2407 218 2412 227
rect 2384 215 2392 218
rect 2378 200 2392 215
rect 2394 205 2402 218
rect 2394 201 2396 205
rect 2400 201 2402 205
rect 2394 200 2402 201
rect 2404 212 2412 218
rect 2404 208 2406 212
rect 2410 208 2412 212
rect 2404 200 2412 208
rect 2414 221 2419 227
rect 2414 220 2421 221
rect 2414 216 2416 220
rect 2420 216 2421 220
rect 2414 215 2421 216
rect 2414 200 2419 215
rect 2455 206 2460 227
rect 2453 205 2460 206
rect 2453 201 2454 205
rect 2458 201 2460 205
rect 2453 200 2460 201
rect 2462 226 2474 227
rect 2462 222 2464 226
rect 2468 222 2474 226
rect 2462 219 2474 222
rect 2462 215 2464 219
rect 2468 218 2474 219
rect 2491 218 2496 227
rect 2468 215 2476 218
rect 2462 200 2476 215
rect 2478 205 2486 218
rect 2478 201 2480 205
rect 2484 201 2486 205
rect 2478 200 2486 201
rect 2488 212 2496 218
rect 2488 208 2490 212
rect 2494 208 2496 212
rect 2488 200 2496 208
rect 2498 221 2503 227
rect 2498 220 2505 221
rect 2498 216 2500 220
rect 2504 216 2505 220
rect 2498 215 2505 216
rect 2498 200 2503 215
rect 2517 205 2522 211
rect 2515 204 2522 205
rect 2515 200 2516 204
rect 2520 200 2522 204
rect 2515 199 2522 200
rect 2524 209 2530 211
rect 2524 204 2532 209
rect 2524 200 2526 204
rect 2530 200 2532 204
rect 2524 199 2532 200
rect 2534 204 2542 209
rect 2534 200 2536 204
rect 2540 200 2542 204
rect 2534 199 2542 200
rect 2544 208 2551 209
rect 2612 208 2617 214
rect 2544 204 2546 208
rect 2550 204 2551 208
rect 2544 199 2551 204
rect 2610 207 2617 208
rect 2610 203 2611 207
rect 2615 203 2617 207
rect 2610 202 2617 203
rect 2619 212 2625 214
rect 2619 207 2627 212
rect 2619 203 2621 207
rect 2625 203 2627 207
rect 2619 202 2627 203
rect 2629 207 2637 212
rect 2629 203 2631 207
rect 2635 203 2637 207
rect 2629 202 2637 203
rect 2639 211 2646 212
rect 2639 207 2641 211
rect 2645 207 2646 211
rect 2698 209 2703 230
rect 2639 202 2646 207
rect 2696 208 2703 209
rect 2696 204 2697 208
rect 2701 204 2703 208
rect 2696 203 2703 204
rect 2705 229 2717 230
rect 2705 225 2707 229
rect 2711 225 2717 229
rect 2705 222 2717 225
rect 2705 218 2707 222
rect 2711 221 2717 222
rect 2734 221 2739 230
rect 2711 218 2719 221
rect 2705 203 2719 218
rect 2721 208 2729 221
rect 2721 204 2723 208
rect 2727 204 2729 208
rect 2721 203 2729 204
rect 2731 215 2739 221
rect 2731 211 2733 215
rect 2737 211 2739 215
rect 2731 203 2739 211
rect 2741 224 2746 230
rect 2741 223 2748 224
rect 2741 219 2743 223
rect 2747 219 2748 223
rect 2741 218 2748 219
rect 2741 203 2746 218
rect 2782 209 2787 230
rect 2780 208 2787 209
rect 2780 204 2781 208
rect 2785 204 2787 208
rect 2780 203 2787 204
rect 2789 229 2801 230
rect 2789 225 2791 229
rect 2795 225 2801 229
rect 2789 222 2801 225
rect 2789 218 2791 222
rect 2795 221 2801 222
rect 2818 221 2823 230
rect 2795 218 2803 221
rect 2789 203 2803 218
rect 2805 208 2813 221
rect 2805 204 2807 208
rect 2811 204 2813 208
rect 2805 203 2813 204
rect 2815 215 2823 221
rect 2815 211 2817 215
rect 2821 211 2823 215
rect 2815 203 2823 211
rect 2825 224 2830 230
rect 2825 223 2832 224
rect 2825 219 2827 223
rect 2831 219 2832 223
rect 2825 218 2832 219
rect 2825 203 2830 218
rect 2844 208 2849 214
rect 2842 207 2849 208
rect 2842 203 2843 207
rect 2847 203 2849 207
rect 2842 202 2849 203
rect 2851 212 2857 214
rect 2851 207 2859 212
rect 2851 203 2853 207
rect 2857 203 2859 207
rect 2851 202 2859 203
rect 2861 207 2869 212
rect 2861 203 2863 207
rect 2867 203 2869 207
rect 2861 202 2869 203
rect 2871 211 2878 212
rect 2871 207 2873 211
rect 2877 207 2878 211
rect 2871 202 2878 207
rect 1794 154 1811 155
rect 1794 150 1795 154
rect 1799 150 1802 154
rect 1806 153 1811 154
rect 1806 150 1819 153
rect 1794 148 1819 150
rect 1794 143 1819 146
rect 592 128 599 136
rect 572 121 578 128
rect 1457 128 1462 135
rect 1455 127 1462 128
rect 1455 123 1456 127
rect 1460 123 1462 127
rect 1455 122 1462 123
rect 1166 120 1181 121
rect 1170 116 1181 120
rect 1166 115 1181 116
rect 1183 120 1203 121
rect 1183 116 1199 120
rect 1183 115 1203 116
rect 1210 120 1220 121
rect 1210 116 1212 120
rect 1216 116 1220 120
rect 1210 115 1220 116
rect 1222 120 1241 121
rect 1222 116 1229 120
rect 1233 116 1241 120
rect 1222 115 1241 116
rect 1243 120 1251 121
rect 1243 116 1246 120
rect 1250 116 1251 120
rect 1243 115 1251 116
rect 1264 120 1274 121
rect 1264 116 1266 120
rect 1270 116 1274 120
rect 1264 115 1274 116
rect 1276 120 1295 121
rect 1276 116 1283 120
rect 1287 116 1295 120
rect 1276 115 1295 116
rect 1297 120 1305 121
rect 1297 116 1300 120
rect 1304 116 1305 120
rect 1297 115 1305 116
rect 1320 120 1330 121
rect 1320 116 1322 120
rect 1326 116 1330 120
rect 1320 115 1330 116
rect 1332 120 1351 121
rect 1332 116 1339 120
rect 1343 116 1351 120
rect 1332 115 1351 116
rect 1353 120 1361 121
rect 1353 116 1356 120
rect 1360 116 1361 120
rect 1353 115 1361 116
rect 1374 120 1384 121
rect 1374 116 1376 120
rect 1380 116 1384 120
rect 1374 115 1384 116
rect 1386 120 1405 121
rect 1386 116 1393 120
rect 1397 116 1405 120
rect 1386 115 1405 116
rect 1407 120 1415 121
rect 1407 116 1410 120
rect 1414 116 1415 120
rect 1457 118 1462 122
rect 1464 118 1474 135
rect 1407 115 1415 116
rect 1466 109 1474 118
rect 1466 105 1467 109
rect 1471 107 1474 109
rect 1476 127 1481 135
rect 1794 139 1815 143
rect 1794 137 1819 139
rect 1794 135 1807 137
rect 1794 131 1807 133
rect 1794 130 1795 131
rect 1476 126 1483 127
rect 1476 122 1478 126
rect 1482 122 1483 126
rect 1476 119 1483 122
rect 1476 115 1478 119
rect 1482 115 1483 119
rect 1791 127 1795 130
rect 1799 130 1807 131
rect 1799 127 1816 130
rect 1791 125 1816 127
rect 1791 118 1816 123
rect 1476 114 1483 115
rect 1476 107 1481 114
rect 1708 109 1718 110
rect 1471 105 1472 107
rect 1466 104 1472 105
rect 1708 105 1709 109
rect 1713 105 1718 109
rect 1708 103 1718 105
rect 1708 99 1718 101
rect 1708 95 1713 99
rect 1717 95 1718 99
rect 1791 114 1816 116
rect 1791 108 1819 114
rect 2066 113 2074 116
rect 2049 108 2054 113
rect 1791 104 1807 108
rect 1811 104 1814 108
rect 1818 104 1819 108
rect 1791 100 1819 104
rect 2047 107 2054 108
rect 2047 103 2048 107
rect 2052 103 2054 107
rect 2047 102 2054 103
rect 1791 96 1819 98
rect 1708 93 1718 95
rect 1791 92 1799 96
rect 1803 92 1806 96
rect 1810 92 1819 96
rect 2049 95 2054 102
rect 2056 95 2061 113
rect 2063 104 2074 113
rect 2076 110 2081 116
rect 2722 118 2730 121
rect 2395 115 2403 118
rect 2378 110 2383 115
rect 2076 109 2083 110
rect 2076 105 2078 109
rect 2082 105 2083 109
rect 2076 104 2083 105
rect 2376 109 2383 110
rect 2376 105 2377 109
rect 2381 105 2383 109
rect 2376 104 2383 105
rect 2063 100 2072 104
rect 2063 96 2066 100
rect 2070 96 2072 100
rect 2063 95 2072 96
rect 2378 97 2383 104
rect 2385 97 2390 115
rect 2392 106 2403 115
rect 2405 112 2410 118
rect 2705 113 2710 118
rect 2703 112 2710 113
rect 2405 111 2412 112
rect 2405 107 2407 111
rect 2411 107 2412 111
rect 2703 108 2704 112
rect 2708 108 2710 112
rect 2703 107 2710 108
rect 2405 106 2412 107
rect 2392 102 2401 106
rect 2392 98 2395 102
rect 2399 98 2401 102
rect 2705 100 2710 107
rect 2712 100 2717 118
rect 2719 109 2730 118
rect 2732 115 2737 121
rect 2732 114 2739 115
rect 2732 110 2734 114
rect 2738 110 2739 114
rect 2732 109 2739 110
rect 2719 105 2728 109
rect 2719 101 2722 105
rect 2726 101 2728 105
rect 2719 100 2728 101
rect 2392 97 2401 98
rect 1708 89 1718 91
rect 1706 85 1713 89
rect 1717 85 1718 89
rect 1706 83 1718 85
rect 1791 90 1819 92
rect 1791 86 1819 88
rect 1791 82 1807 86
rect 1811 82 1814 86
rect 1818 82 1819 86
rect 1706 79 1718 81
rect 1706 76 1713 79
rect 1712 75 1713 76
rect 1717 75 1718 79
rect 1712 74 1718 75
rect 1791 80 1819 82
rect 1791 76 1819 78
rect 1791 72 1792 76
rect 1796 72 1799 76
rect 1803 73 1819 76
rect 1803 72 1804 73
rect 1791 71 1804 72
rect 2259 68 2265 70
rect 2250 63 2255 68
rect 2248 62 2255 63
rect 2248 58 2249 62
rect 2253 58 2255 62
rect 2248 55 2255 58
rect 2248 51 2249 55
rect 2253 51 2255 55
rect 2248 50 2255 51
rect 2257 67 2265 68
rect 2257 63 2259 67
rect 2263 63 2265 67
rect 2257 57 2265 63
rect 2267 69 2275 70
rect 2267 65 2269 69
rect 2273 65 2275 69
rect 2267 62 2275 65
rect 2267 58 2269 62
rect 2273 58 2275 62
rect 2267 57 2275 58
rect 2277 69 2284 70
rect 2277 65 2279 69
rect 2283 65 2284 69
rect 2352 68 2358 70
rect 2277 57 2284 65
rect 2343 63 2348 68
rect 2341 62 2348 63
rect 2341 58 2342 62
rect 2346 58 2348 62
rect 2257 50 2263 57
rect 2341 55 2348 58
rect 2341 51 2342 55
rect 2346 51 2348 55
rect 2341 50 2348 51
rect 2350 67 2358 68
rect 2350 63 2352 67
rect 2356 63 2358 67
rect 2350 57 2358 63
rect 2360 69 2368 70
rect 2360 65 2362 69
rect 2366 65 2368 69
rect 2360 62 2368 65
rect 2360 58 2362 62
rect 2366 58 2368 62
rect 2360 57 2368 58
rect 2370 69 2377 70
rect 2370 65 2372 69
rect 2376 65 2377 69
rect 2439 68 2445 70
rect 2370 57 2377 65
rect 2430 63 2435 68
rect 2428 62 2435 63
rect 2428 58 2429 62
rect 2433 58 2435 62
rect 2350 50 2356 57
rect 2428 55 2435 58
rect 2428 51 2429 55
rect 2433 51 2435 55
rect 2428 50 2435 51
rect 2437 67 2445 68
rect 2437 63 2439 67
rect 2443 63 2445 67
rect 2437 57 2445 63
rect 2447 69 2455 70
rect 2447 65 2449 69
rect 2453 65 2455 69
rect 2447 62 2455 65
rect 2447 58 2449 62
rect 2453 58 2455 62
rect 2447 57 2455 58
rect 2457 69 2464 70
rect 2457 65 2459 69
rect 2463 65 2464 69
rect 2457 57 2464 65
rect 2437 50 2443 57
<< metal1 >>
rect 1549 1139 1554 1140
rect 1549 1133 1957 1139
rect 1549 1107 1554 1133
rect 1817 1105 1912 1110
rect 1858 1097 1921 1100
rect 1600 1090 1803 1093
rect 1601 1080 1605 1090
rect 1539 1063 1563 1064
rect 1539 1062 1692 1063
rect 1539 1059 1698 1062
rect 76 1042 517 1046
rect 76 1020 80 1042
rect 559 1040 821 1044
rect 158 1033 159 1036
rect 559 1038 563 1040
rect 510 1035 563 1038
rect 374 1033 500 1034
rect 573 1033 617 1035
rect 158 1032 500 1033
rect 153 1031 500 1032
rect 567 1032 617 1033
rect 666 1032 710 1035
rect 753 1034 797 1035
rect 753 1032 805 1034
rect 567 1031 805 1032
rect 153 1029 579 1031
rect 153 1025 177 1029
rect 181 1025 187 1029
rect 191 1025 264 1029
rect 268 1025 274 1029
rect 278 1025 357 1029
rect 361 1025 367 1029
rect 371 1028 579 1029
rect 371 1025 377 1028
rect 573 1027 579 1028
rect 583 1027 589 1031
rect 593 1028 672 1031
rect 593 1027 617 1028
rect 666 1027 672 1028
rect 676 1027 682 1031
rect 686 1028 759 1031
rect 686 1027 710 1028
rect 753 1027 759 1028
rect 763 1027 769 1031
rect 773 1028 805 1031
rect 773 1027 797 1028
rect 817 1025 821 1040
rect 994 1036 1409 1039
rect 994 1035 1045 1036
rect 1037 1025 1042 1028
rect 510 1020 541 1024
rect 157 1015 158 1019
rect 162 1015 177 1019
rect 157 1008 169 1012
rect 164 1003 169 1008
rect 173 1011 177 1015
rect 181 1017 193 1020
rect 181 1014 188 1017
rect 192 1013 193 1017
rect 244 1015 245 1019
rect 249 1015 264 1019
rect 188 1012 193 1013
rect 173 1007 185 1011
rect 181 1003 185 1007
rect 164 999 171 1003
rect 175 999 178 1003
rect 157 986 161 995
rect 165 991 170 995
rect 181 988 185 999
rect 189 998 193 1012
rect 245 1008 256 1012
rect 251 1003 256 1008
rect 260 1011 264 1015
rect 268 1017 280 1020
rect 268 1014 275 1017
rect 279 1013 280 1017
rect 337 1015 338 1019
rect 342 1015 357 1019
rect 275 1012 280 1013
rect 260 1007 272 1011
rect 268 1003 272 1007
rect 251 999 258 1003
rect 262 999 265 1003
rect 189 995 218 998
rect 189 994 193 995
rect 150 982 161 986
rect 168 986 185 988
rect 172 984 185 986
rect 188 993 193 994
rect 192 989 193 993
rect 188 986 193 989
rect 168 979 172 982
rect 192 982 193 986
rect 188 981 193 982
rect 157 975 158 979
rect 162 975 163 979
rect 157 969 163 975
rect 168 974 172 975
rect 177 977 178 981
rect 182 977 183 981
rect 177 969 183 977
rect 153 965 187 969
rect 191 965 197 969
rect 153 961 197 965
rect 154 954 158 961
rect 214 959 218 995
rect 244 985 248 995
rect 252 991 257 995
rect 268 988 272 999
rect 276 994 280 1012
rect 338 1008 349 1012
rect 344 1003 349 1008
rect 353 1011 357 1015
rect 361 1017 373 1020
rect 577 1019 589 1022
rect 361 1014 368 1017
rect 372 1013 373 1017
rect 386 1013 558 1017
rect 563 1013 564 1017
rect 577 1015 578 1019
rect 582 1016 589 1019
rect 593 1017 608 1021
rect 612 1017 613 1021
rect 670 1019 682 1022
rect 577 1014 582 1015
rect 368 1012 373 1013
rect 353 1007 365 1011
rect 361 1003 365 1007
rect 344 999 351 1003
rect 355 999 358 1003
rect 241 982 248 985
rect 255 986 272 988
rect 259 984 272 986
rect 275 993 280 994
rect 279 989 280 993
rect 275 986 280 989
rect 255 979 259 982
rect 279 984 280 986
rect 279 982 286 984
rect 275 981 286 982
rect 337 985 341 995
rect 345 991 350 995
rect 361 988 365 999
rect 369 1005 373 1012
rect 577 1007 581 1014
rect 593 1013 597 1017
rect 670 1015 671 1019
rect 675 1016 682 1019
rect 686 1017 701 1021
rect 705 1017 706 1021
rect 757 1019 769 1022
rect 817 1021 1023 1025
rect 670 1014 675 1015
rect 369 1001 455 1005
rect 521 1003 581 1007
rect 369 994 373 1001
rect 577 996 581 1003
rect 585 1009 597 1013
rect 601 1011 612 1014
rect 585 1005 589 1009
rect 601 1005 606 1011
rect 592 1001 595 1005
rect 599 1001 606 1005
rect 670 1003 674 1014
rect 686 1013 690 1017
rect 757 1015 758 1019
rect 762 1016 769 1019
rect 773 1017 788 1021
rect 792 1017 793 1021
rect 757 1014 762 1015
rect 577 995 582 996
rect 334 982 341 985
rect 348 986 365 988
rect 352 984 365 986
rect 368 993 373 994
rect 372 989 373 993
rect 386 991 559 994
rect 577 991 578 995
rect 368 986 373 989
rect 244 975 245 979
rect 249 975 250 979
rect 244 969 250 975
rect 255 974 259 975
rect 264 977 265 981
rect 269 977 270 981
rect 348 979 352 982
rect 372 982 373 986
rect 577 988 582 991
rect 577 984 578 988
rect 585 990 589 1001
rect 647 1000 674 1003
rect 600 993 605 997
rect 585 988 602 990
rect 585 986 598 988
rect 577 983 582 984
rect 609 987 613 997
rect 647 988 651 1000
rect 609 984 616 987
rect 368 981 373 982
rect 264 969 270 977
rect 337 975 338 979
rect 342 975 343 979
rect 337 969 343 975
rect 348 974 352 975
rect 357 977 358 981
rect 362 977 363 981
rect 587 979 588 983
rect 592 979 593 983
rect 357 969 363 977
rect 386 973 560 976
rect 587 971 593 979
rect 598 981 602 984
rect 670 996 674 1000
rect 678 1009 690 1013
rect 694 1013 708 1014
rect 694 1011 705 1013
rect 678 1005 682 1009
rect 694 1005 699 1011
rect 685 1001 688 1005
rect 692 1001 699 1005
rect 670 995 675 996
rect 670 991 671 995
rect 670 988 675 991
rect 670 984 671 988
rect 678 990 682 1001
rect 757 1000 761 1014
rect 773 1013 777 1017
rect 693 993 698 997
rect 678 988 695 990
rect 678 986 691 988
rect 670 983 675 984
rect 702 987 706 997
rect 735 996 761 1000
rect 765 1009 777 1013
rect 781 1013 795 1014
rect 1037 1013 1040 1025
rect 1059 1017 1062 1036
rect 1072 1025 1126 1028
rect 1104 1019 1108 1021
rect 781 1011 792 1013
rect 765 1005 769 1009
rect 781 1005 786 1011
rect 796 1009 1041 1013
rect 772 1001 775 1005
rect 779 1001 786 1005
rect 1104 1002 1108 1013
rect 1123 1010 1126 1025
rect 1142 1017 1145 1036
rect 1205 1017 1208 1036
rect 1215 1031 1218 1036
rect 1259 1017 1262 1036
rect 1269 1031 1272 1036
rect 1315 1017 1318 1036
rect 1325 1031 1328 1036
rect 1369 1017 1372 1036
rect 1379 1031 1382 1036
rect 1123 1007 1173 1010
rect 702 984 709 987
rect 721 986 722 990
rect 598 976 602 977
rect 607 977 608 981
rect 612 977 613 981
rect 607 971 613 977
rect 680 979 681 983
rect 685 979 686 983
rect 680 971 686 979
rect 691 981 695 984
rect 691 976 695 977
rect 700 977 701 981
rect 705 977 706 981
rect 700 971 706 977
rect 240 965 274 969
rect 278 965 284 969
rect 240 964 284 965
rect 333 965 367 969
rect 371 965 377 969
rect 240 961 267 964
rect 333 961 377 965
rect 573 967 579 971
rect 583 967 617 971
rect 666 967 672 971
rect 676 967 710 971
rect 573 963 617 967
rect 242 954 246 961
rect 279 957 312 960
rect 333 954 337 961
rect 609 959 613 963
rect 628 962 658 965
rect 666 963 710 967
rect 721 966 725 986
rect 567 958 671 959
rect 567 956 693 958
rect 702 956 706 963
rect 735 965 739 996
rect 757 995 762 996
rect 757 991 758 995
rect 745 966 749 986
rect 757 988 762 991
rect 757 984 758 988
rect 765 990 769 1001
rect 780 993 785 997
rect 765 988 782 990
rect 765 986 778 988
rect 757 983 762 984
rect 789 988 793 997
rect 1087 998 1090 1001
rect 1104 992 1107 1002
rect 1159 997 1162 1000
rect 789 984 797 988
rect 767 979 768 983
rect 772 979 773 983
rect 767 971 773 979
rect 778 981 782 984
rect 778 976 782 977
rect 787 977 788 981
rect 792 977 793 981
rect 787 971 793 977
rect 753 967 759 971
rect 763 967 797 971
rect 753 963 797 967
rect 791 956 795 963
rect 988 959 992 992
rect 1104 988 1105 992
rect 1104 980 1107 988
rect 1169 987 1173 1007
rect 1176 991 1179 1013
rect 1189 1008 1192 1013
rect 1222 1008 1225 1013
rect 1189 1005 1225 1008
rect 1191 997 1193 1000
rect 1205 998 1209 1000
rect 1213 998 1214 1000
rect 1205 997 1214 998
rect 1176 987 1177 991
rect 1205 989 1208 997
rect 1222 996 1225 1005
rect 1243 1008 1246 1013
rect 1276 1008 1279 1013
rect 1243 1005 1279 1008
rect 1299 1008 1302 1013
rect 1332 1008 1335 1013
rect 1299 1005 1335 1008
rect 1353 1008 1356 1013
rect 1386 1008 1389 1013
rect 1353 1005 1389 1008
rect 1229 996 1232 1005
rect 1243 1000 1250 1001
rect 1243 998 1247 1000
rect 1264 996 1268 999
rect 1222 993 1232 996
rect 1205 987 1210 989
rect 1176 979 1179 987
rect 1205 986 1206 987
rect 1222 980 1225 993
rect 1264 992 1267 996
rect 1276 993 1279 1005
rect 1332 1004 1335 1005
rect 1300 997 1303 1000
rect 1276 990 1295 993
rect 1276 980 1279 990
rect 1324 994 1327 996
rect 1312 986 1315 992
rect 1326 990 1327 994
rect 1324 989 1327 990
rect 1289 983 1315 986
rect 1332 980 1335 1000
rect 1356 996 1357 999
rect 1375 1000 1381 1001
rect 1375 998 1378 1000
rect 1356 987 1359 996
rect 1386 995 1389 1005
rect 1358 983 1359 987
rect 1386 980 1389 991
rect 1070 970 1073 976
rect 1142 970 1145 975
rect 1188 970 1191 976
rect 1242 970 1245 976
rect 1298 970 1301 976
rect 1352 970 1355 976
rect 1046 967 1391 970
rect 805 956 1007 959
rect 349 955 1007 956
rect 349 954 737 955
rect 45 953 272 954
rect 285 953 737 954
rect 45 952 737 953
rect 45 950 410 952
rect 45 946 81 950
rect 85 946 95 950
rect 99 946 109 950
rect 113 947 192 950
rect 113 946 176 947
rect 45 835 49 946
rect 65 945 80 946
rect 79 926 83 933
rect 79 925 84 926
rect 79 921 80 925
rect 87 925 91 946
rect 94 940 107 941
rect 94 936 97 940
rect 101 936 103 940
rect 94 935 107 936
rect 94 928 100 935
rect 110 929 114 946
rect 180 946 192 947
rect 196 947 276 950
rect 196 946 260 947
rect 157 935 169 941
rect 176 940 180 943
rect 264 946 276 947
rect 280 946 313 950
rect 317 946 327 950
rect 331 946 341 950
rect 345 948 410 950
rect 414 948 424 952
rect 428 948 438 952
rect 442 949 521 952
rect 442 948 505 949
rect 345 946 380 948
rect 190 937 212 941
rect 216 937 217 941
rect 241 940 253 941
rect 190 936 194 937
rect 176 935 180 936
rect 157 932 162 935
rect 157 931 158 932
rect 87 921 90 925
rect 94 921 95 925
rect 99 921 100 925
rect 104 921 105 925
rect 110 924 114 925
rect 149 928 158 931
rect 183 932 194 936
rect 241 936 246 940
rect 250 936 253 940
rect 241 935 253 936
rect 260 940 264 943
rect 274 937 296 941
rect 300 937 301 941
rect 274 936 278 937
rect 260 935 264 936
rect 183 928 187 932
rect 201 929 202 933
rect 206 929 217 933
rect 79 920 84 921
rect 79 912 83 920
rect 99 916 105 921
rect 86 912 87 916
rect 91 912 105 916
rect 111 914 115 917
rect 149 914 152 928
rect 157 927 162 928
rect 166 926 187 928
rect 79 903 83 908
rect 79 902 84 903
rect 79 898 80 902
rect 84 898 91 901
rect 79 895 91 898
rect 95 899 99 912
rect 158 922 166 923
rect 170 924 187 926
rect 158 919 170 922
rect 111 908 115 910
rect 102 904 106 908
rect 110 904 115 908
rect 102 903 115 904
rect 158 907 162 919
rect 183 917 187 924
rect 191 922 192 926
rect 196 925 197 926
rect 196 922 208 925
rect 191 921 208 922
rect 204 918 208 921
rect 204 917 209 918
rect 172 911 178 916
rect 183 913 195 917
rect 199 913 200 917
rect 204 913 205 917
rect 172 909 174 911
rect 165 907 174 909
rect 204 912 209 913
rect 213 913 217 929
rect 241 932 246 935
rect 241 928 242 932
rect 267 932 278 936
rect 267 928 271 932
rect 285 929 286 933
rect 290 930 301 933
rect 290 929 304 930
rect 241 927 246 928
rect 250 926 271 928
rect 297 927 304 929
rect 242 922 250 923
rect 254 924 271 926
rect 242 919 254 922
rect 204 908 208 912
rect 165 903 178 907
rect 184 904 208 908
rect 213 909 215 913
rect 158 902 162 903
rect 184 902 188 904
rect 95 895 109 899
rect 113 895 114 899
rect 171 895 172 899
rect 176 895 177 899
rect 213 900 217 909
rect 242 907 246 919
rect 267 917 271 924
rect 275 922 276 926
rect 280 925 281 926
rect 280 922 292 925
rect 275 921 292 922
rect 288 918 292 921
rect 288 917 293 918
rect 256 911 262 916
rect 267 913 279 917
rect 283 913 284 917
rect 288 913 289 917
rect 256 909 258 911
rect 249 907 258 909
rect 288 912 293 913
rect 288 908 292 912
rect 249 903 262 907
rect 268 904 292 908
rect 242 902 246 903
rect 268 902 272 904
rect 184 897 188 898
rect 193 896 194 900
rect 198 896 217 900
rect 171 890 177 895
rect 255 895 256 899
rect 260 895 261 899
rect 297 900 301 927
rect 311 926 315 933
rect 311 925 316 926
rect 311 921 312 925
rect 319 925 323 946
rect 326 940 339 941
rect 326 936 329 940
rect 333 936 335 940
rect 326 935 339 936
rect 326 928 332 935
rect 342 929 346 946
rect 354 927 365 930
rect 319 921 322 925
rect 326 921 327 925
rect 331 921 332 925
rect 336 921 337 925
rect 342 924 346 925
rect 311 920 316 921
rect 311 912 315 920
rect 331 916 337 921
rect 318 912 319 916
rect 323 912 337 916
rect 343 915 347 917
rect 268 897 272 898
rect 277 896 278 900
rect 282 896 301 900
rect 305 909 315 912
rect 305 897 308 909
rect 255 890 261 895
rect 311 903 315 909
rect 311 902 316 903
rect 311 898 312 902
rect 316 898 323 901
rect 311 895 323 898
rect 327 899 331 912
rect 343 908 347 911
rect 334 904 338 908
rect 342 904 347 908
rect 334 903 347 904
rect 327 895 341 899
rect 345 895 346 899
rect 78 886 81 890
rect 85 886 91 890
rect 95 886 159 890
rect 163 886 212 890
rect 216 886 243 890
rect 247 886 296 890
rect 300 886 313 890
rect 317 886 323 890
rect 327 889 351 890
rect 327 886 345 889
rect 64 883 345 886
rect 64 882 351 883
rect 168 880 212 882
rect 168 876 174 880
rect 178 876 202 880
rect 206 876 212 880
rect 172 868 178 876
rect 172 864 173 868
rect 177 864 178 868
rect 183 868 187 869
rect 192 868 198 876
rect 192 864 193 868
rect 197 864 198 868
rect 203 868 208 871
rect 207 864 208 868
rect 183 861 187 864
rect 203 863 208 864
rect 183 857 200 861
rect 172 845 176 855
rect 180 850 185 854
rect 196 853 200 857
rect 180 842 186 846
rect 190 842 193 846
rect 44 815 49 835
rect 180 836 184 842
rect 196 838 200 849
rect 167 833 184 836
rect 188 834 200 838
rect 204 859 365 863
rect 188 830 192 834
rect 204 833 208 859
rect 374 837 378 946
rect 408 928 412 935
rect 408 927 413 928
rect 408 923 409 927
rect 416 927 420 948
rect 423 942 436 943
rect 423 938 426 942
rect 430 938 432 942
rect 423 937 436 938
rect 423 930 429 937
rect 439 931 443 948
rect 509 948 521 949
rect 525 949 605 952
rect 525 948 589 949
rect 486 937 498 943
rect 505 942 509 945
rect 593 948 605 949
rect 609 948 642 952
rect 646 948 656 952
rect 660 948 670 952
rect 674 951 737 952
rect 741 951 751 955
rect 755 951 765 955
rect 769 952 848 955
rect 769 951 832 952
rect 674 948 710 951
rect 519 939 541 943
rect 545 939 546 943
rect 561 942 582 943
rect 519 938 523 939
rect 505 937 509 938
rect 486 934 491 937
rect 416 923 419 927
rect 423 923 424 927
rect 428 923 429 927
rect 433 923 434 927
rect 439 926 443 927
rect 486 933 487 934
rect 408 922 413 923
rect 408 914 412 922
rect 428 918 434 923
rect 415 914 416 918
rect 420 914 434 918
rect 440 916 444 919
rect 408 905 412 910
rect 408 904 413 905
rect 408 900 409 904
rect 413 900 420 903
rect 408 897 420 900
rect 424 901 428 914
rect 440 910 444 912
rect 431 906 435 910
rect 439 906 444 910
rect 431 905 444 906
rect 424 897 438 901
rect 442 897 443 901
rect 461 901 465 929
rect 478 930 487 933
rect 512 934 523 938
rect 561 938 575 942
rect 579 938 582 942
rect 561 937 582 938
rect 589 942 593 945
rect 603 939 625 943
rect 629 939 630 943
rect 603 938 607 939
rect 589 937 593 938
rect 512 930 516 934
rect 530 931 531 935
rect 535 931 546 935
rect 478 916 481 930
rect 486 929 491 930
rect 495 928 516 930
rect 487 924 495 925
rect 499 926 516 928
rect 487 921 499 924
rect 487 909 491 921
rect 512 919 516 926
rect 520 924 521 928
rect 525 927 526 928
rect 525 924 537 927
rect 520 923 537 924
rect 533 920 537 923
rect 533 919 538 920
rect 501 913 507 918
rect 512 915 524 919
rect 528 915 529 919
rect 533 915 534 919
rect 501 911 503 913
rect 494 909 503 911
rect 533 914 538 915
rect 542 915 546 931
rect 570 934 575 937
rect 570 930 571 934
rect 596 934 607 938
rect 596 930 600 934
rect 614 931 615 935
rect 619 931 632 935
rect 570 929 575 930
rect 579 928 600 930
rect 571 924 579 925
rect 583 926 600 928
rect 571 921 583 924
rect 533 910 537 914
rect 494 905 507 909
rect 513 906 537 910
rect 542 911 544 915
rect 487 904 491 905
rect 513 904 517 906
rect 457 898 465 901
rect 500 897 501 901
rect 505 897 506 901
rect 542 902 546 911
rect 571 909 575 921
rect 596 919 600 926
rect 604 924 605 928
rect 609 927 610 928
rect 609 924 621 927
rect 604 923 621 924
rect 617 920 621 923
rect 617 919 622 920
rect 585 913 591 918
rect 596 915 608 919
rect 612 915 613 919
rect 617 915 618 919
rect 585 911 587 913
rect 578 909 587 911
rect 617 914 622 915
rect 617 910 621 914
rect 578 905 591 909
rect 597 906 621 910
rect 571 904 575 905
rect 597 904 601 906
rect 513 899 517 900
rect 522 898 523 902
rect 527 898 546 902
rect 500 892 506 897
rect 584 897 585 901
rect 589 897 590 901
rect 626 902 630 931
rect 640 928 644 935
rect 640 927 645 928
rect 640 923 641 927
rect 648 927 652 948
rect 655 942 668 943
rect 655 938 658 942
rect 662 938 664 942
rect 655 937 668 938
rect 655 930 661 937
rect 671 931 675 948
rect 648 923 651 927
rect 655 923 656 927
rect 660 923 661 927
rect 665 923 666 927
rect 671 926 675 927
rect 640 922 645 923
rect 640 914 644 922
rect 660 918 666 923
rect 647 914 648 918
rect 652 914 666 918
rect 672 917 676 919
rect 597 899 601 900
rect 606 898 607 902
rect 611 898 630 902
rect 634 911 644 914
rect 634 899 637 911
rect 584 892 590 897
rect 640 905 644 911
rect 640 904 645 905
rect 640 900 641 904
rect 645 900 652 903
rect 640 897 652 900
rect 656 901 660 914
rect 672 910 676 913
rect 663 906 667 910
rect 671 906 676 910
rect 663 905 676 906
rect 656 897 670 901
rect 674 897 675 901
rect 407 888 410 892
rect 414 888 420 892
rect 424 888 488 892
rect 492 888 541 892
rect 545 888 572 892
rect 576 888 625 892
rect 629 888 642 892
rect 646 888 652 892
rect 656 891 680 892
rect 656 888 672 891
rect 407 887 672 888
rect 392 885 672 887
rect 678 885 680 891
rect 392 884 680 885
rect 392 883 408 884
rect 497 882 541 884
rect 497 878 503 882
rect 507 878 531 882
rect 535 878 541 882
rect 501 870 507 878
rect 501 866 502 870
rect 506 866 507 870
rect 512 870 516 871
rect 521 870 527 878
rect 521 866 522 870
rect 526 866 527 870
rect 532 870 537 873
rect 627 871 698 874
rect 536 866 537 870
rect 512 863 516 866
rect 532 865 537 866
rect 394 859 462 863
rect 512 859 529 863
rect 501 847 505 857
rect 509 852 514 856
rect 525 855 529 859
rect 509 844 515 848
rect 519 844 522 848
rect 203 832 208 833
rect 172 826 173 830
rect 177 826 192 830
rect 195 828 203 830
rect 207 828 208 832
rect 195 826 208 828
rect 190 820 191 823
rect 168 819 191 820
rect 195 820 196 823
rect 195 819 202 820
rect 168 816 202 819
rect 206 816 212 820
rect 168 815 212 816
rect 373 817 378 837
rect 509 838 513 844
rect 525 840 529 851
rect 496 835 513 838
rect 517 836 529 840
rect 533 859 537 865
rect 533 856 684 859
rect 688 856 689 859
rect 517 832 521 836
rect 533 835 537 856
rect 532 834 537 835
rect 501 828 502 832
rect 506 828 521 832
rect 524 830 532 832
rect 536 830 537 834
rect 524 828 537 830
rect 519 822 520 825
rect 497 821 520 822
rect 524 822 525 825
rect 524 821 531 822
rect 497 818 531 821
rect 535 818 541 822
rect 497 817 541 818
rect 44 812 212 815
rect 44 811 172 812
rect 350 811 365 815
rect 169 808 172 811
rect 373 814 541 817
rect 373 813 499 814
rect 496 810 499 813
rect 44 804 350 808
rect 44 800 80 804
rect 84 800 94 804
rect 98 800 108 804
rect 112 801 191 804
rect 112 800 175 801
rect 44 689 48 800
rect 78 780 82 787
rect 78 779 83 780
rect 78 775 79 779
rect 86 779 90 800
rect 93 794 106 795
rect 93 790 96 794
rect 100 790 102 794
rect 93 789 106 790
rect 93 782 99 789
rect 109 783 113 800
rect 179 800 191 801
rect 195 801 275 804
rect 195 800 259 801
rect 156 789 168 795
rect 175 794 179 797
rect 263 800 275 801
rect 279 800 312 804
rect 316 800 326 804
rect 330 800 340 804
rect 344 800 350 804
rect 373 806 679 810
rect 694 809 697 871
rect 701 840 705 948
rect 735 931 739 938
rect 735 930 740 931
rect 735 926 736 930
rect 743 930 747 951
rect 750 945 763 946
rect 750 941 753 945
rect 757 941 759 945
rect 750 940 763 941
rect 750 933 756 940
rect 766 934 770 951
rect 836 951 848 952
rect 852 952 932 955
rect 852 951 916 952
rect 813 940 825 946
rect 832 945 836 948
rect 920 951 932 952
rect 936 951 969 955
rect 973 951 983 955
rect 987 951 997 955
rect 1001 951 1007 955
rect 846 942 868 946
rect 872 942 873 946
rect 886 945 909 946
rect 846 941 850 942
rect 886 941 902 945
rect 906 941 909 945
rect 832 940 836 941
rect 813 937 818 940
rect 813 936 814 937
rect 743 926 746 930
rect 750 926 751 930
rect 755 926 756 930
rect 760 926 761 930
rect 766 929 770 930
rect 735 925 740 926
rect 735 917 739 925
rect 755 921 761 926
rect 742 917 743 921
rect 747 917 761 921
rect 767 919 771 922
rect 735 908 739 913
rect 735 907 740 908
rect 735 903 736 907
rect 740 903 747 906
rect 735 900 747 903
rect 751 904 755 917
rect 767 913 771 915
rect 758 909 762 913
rect 766 909 771 913
rect 758 908 771 909
rect 751 900 765 904
rect 769 900 770 904
rect 794 902 798 931
rect 805 933 814 936
rect 839 937 850 941
rect 839 933 843 937
rect 857 934 858 938
rect 862 934 873 938
rect 805 919 808 933
rect 813 932 818 933
rect 822 931 843 933
rect 814 927 822 928
rect 826 929 843 931
rect 814 924 826 927
rect 814 912 818 924
rect 839 922 843 929
rect 847 927 848 931
rect 852 930 853 931
rect 852 927 864 930
rect 847 926 864 927
rect 860 923 864 926
rect 860 922 865 923
rect 828 916 834 921
rect 839 918 851 922
rect 855 918 856 922
rect 860 918 861 922
rect 828 914 830 916
rect 821 912 830 914
rect 860 917 865 918
rect 869 918 873 934
rect 860 913 864 917
rect 821 908 834 912
rect 840 909 864 913
rect 869 914 871 918
rect 814 907 818 908
rect 840 907 844 909
rect 794 898 795 902
rect 827 900 828 904
rect 832 900 833 904
rect 869 905 873 914
rect 840 902 844 903
rect 849 901 850 905
rect 854 901 873 905
rect 880 902 883 933
rect 827 895 833 900
rect 887 895 891 941
rect 897 940 909 941
rect 916 945 920 948
rect 930 942 952 946
rect 956 942 957 946
rect 930 941 934 942
rect 916 940 920 941
rect 897 937 902 940
rect 897 933 898 937
rect 923 937 934 941
rect 923 933 927 937
rect 941 934 942 938
rect 946 934 957 938
rect 897 932 902 933
rect 906 931 927 933
rect 898 927 906 928
rect 910 929 927 931
rect 898 924 910 927
rect 898 912 902 924
rect 923 922 927 929
rect 931 927 932 931
rect 936 930 937 931
rect 936 927 948 930
rect 931 926 948 927
rect 944 923 948 926
rect 944 922 949 923
rect 912 916 918 921
rect 923 918 935 922
rect 939 918 940 922
rect 944 918 945 922
rect 912 914 914 916
rect 905 912 914 914
rect 944 917 949 918
rect 944 913 948 917
rect 905 908 918 912
rect 924 909 948 913
rect 898 907 902 908
rect 924 907 928 909
rect 911 900 912 904
rect 916 900 917 904
rect 953 905 957 934
rect 967 931 971 938
rect 967 930 972 931
rect 967 926 968 930
rect 975 930 979 951
rect 982 945 995 946
rect 982 941 985 945
rect 989 941 991 945
rect 982 940 995 941
rect 982 933 988 940
rect 998 934 1002 951
rect 975 926 978 930
rect 982 926 983 930
rect 987 926 988 930
rect 992 926 993 930
rect 998 929 1002 930
rect 967 925 972 926
rect 967 917 971 925
rect 987 921 993 926
rect 974 917 975 921
rect 979 917 993 921
rect 999 920 1003 922
rect 924 902 928 903
rect 933 901 934 905
rect 938 901 957 905
rect 961 914 971 917
rect 961 902 964 914
rect 911 895 917 900
rect 967 908 971 914
rect 967 907 972 908
rect 967 903 968 907
rect 972 903 979 906
rect 967 900 979 903
rect 983 904 987 917
rect 999 913 1003 916
rect 1046 914 1050 967
rect 1214 964 1219 967
rect 1320 964 1324 967
rect 1146 961 1395 964
rect 1146 956 1149 961
rect 1192 955 1195 961
rect 1246 955 1249 961
rect 1302 955 1305 961
rect 1356 955 1359 961
rect 1180 944 1183 952
rect 1180 940 1181 944
rect 990 909 994 913
rect 998 909 1003 913
rect 990 908 1003 909
rect 1014 910 1050 914
rect 983 900 997 904
rect 1001 900 1002 904
rect 734 894 737 895
rect 732 891 737 894
rect 741 891 747 895
rect 751 891 815 895
rect 819 891 868 895
rect 872 891 899 895
rect 903 891 952 895
rect 956 891 969 895
rect 973 891 979 895
rect 983 891 1007 895
rect 1014 891 1018 910
rect 732 889 1018 891
rect 719 887 1018 889
rect 719 886 736 887
rect 719 885 735 886
rect 824 885 868 887
rect 824 881 830 885
rect 834 881 858 885
rect 862 881 868 885
rect 828 873 834 881
rect 828 869 829 873
rect 833 869 834 873
rect 839 873 843 874
rect 848 873 854 881
rect 848 869 849 873
rect 853 869 854 873
rect 859 873 864 876
rect 863 869 864 873
rect 720 856 787 859
rect 791 856 792 859
rect 700 820 705 840
rect 797 828 801 868
rect 839 866 843 869
rect 859 868 864 869
rect 839 862 856 866
rect 809 834 812 861
rect 828 850 832 860
rect 836 855 841 859
rect 852 858 856 862
rect 836 847 842 851
rect 846 847 849 851
rect 836 841 840 847
rect 852 843 856 854
rect 823 838 840 841
rect 844 839 856 843
rect 860 864 864 868
rect 860 861 872 864
rect 844 835 848 839
rect 860 838 864 861
rect 880 840 883 855
rect 859 837 864 838
rect 828 831 829 835
rect 833 831 848 835
rect 851 833 859 835
rect 863 833 864 837
rect 851 831 864 833
rect 846 825 847 828
rect 797 823 801 824
rect 824 824 847 825
rect 851 825 852 828
rect 879 827 884 840
rect 851 824 858 825
rect 824 821 858 824
rect 862 821 868 825
rect 824 820 868 821
rect 1030 825 1033 910
rect 1129 906 1133 934
rect 1163 931 1166 934
rect 1180 918 1183 940
rect 1226 938 1229 951
rect 1226 935 1236 938
rect 1268 935 1271 939
rect 1280 941 1283 951
rect 1280 938 1299 941
rect 1328 941 1331 942
rect 1195 931 1197 934
rect 1217 931 1218 934
rect 1226 926 1229 935
rect 1193 923 1229 926
rect 1193 918 1196 923
rect 1226 918 1229 923
rect 1233 926 1236 935
rect 1247 931 1251 933
rect 1268 932 1272 935
rect 1247 930 1254 931
rect 1280 926 1283 938
rect 1330 937 1331 941
rect 1328 935 1331 937
rect 1304 931 1307 934
rect 1336 931 1339 951
rect 1362 944 1363 948
rect 1360 935 1363 944
rect 1390 940 1393 951
rect 1360 932 1361 935
rect 1379 931 1382 933
rect 1379 930 1385 931
rect 1336 926 1339 927
rect 1390 926 1393 936
rect 1247 923 1283 926
rect 1247 918 1250 923
rect 1280 918 1283 923
rect 1303 923 1339 926
rect 1303 918 1306 923
rect 1336 918 1339 923
rect 1357 923 1393 926
rect 1357 918 1360 923
rect 1390 918 1393 923
rect 1132 904 1133 906
rect 1146 895 1149 914
rect 1209 895 1212 914
rect 1219 895 1222 900
rect 1263 895 1266 914
rect 1273 895 1276 900
rect 1319 895 1322 914
rect 1329 895 1332 900
rect 1373 895 1376 914
rect 1383 895 1386 900
rect 1404 895 1409 1036
rect 1539 940 1543 1059
rect 1674 1057 1698 1059
rect 1674 1056 1715 1057
rect 1674 1052 1694 1056
rect 1698 1053 1715 1056
rect 1719 1053 1720 1057
rect 1727 1054 1729 1058
rect 1733 1054 1741 1058
rect 1736 1053 1741 1054
rect 1603 955 1606 1047
rect 1674 1042 1698 1052
rect 1674 1038 1694 1042
rect 1674 1034 1698 1038
rect 1703 1046 1704 1050
rect 1708 1046 1709 1050
rect 1740 1049 1741 1053
rect 1703 1044 1709 1046
rect 1703 1040 1704 1044
rect 1708 1043 1709 1044
rect 1719 1047 1732 1048
rect 1723 1043 1732 1047
rect 1736 1045 1741 1049
rect 1745 1056 1749 1057
rect 1708 1040 1716 1043
rect 1719 1042 1732 1043
rect 1745 1042 1749 1052
rect 1703 1037 1716 1040
rect 1728 1038 1749 1042
rect 1754 1038 1762 1062
rect 1719 1037 1723 1038
rect 1674 1033 1719 1034
rect 1674 1030 1723 1033
rect 1728 1034 1732 1038
rect 1758 1034 1762 1038
rect 1610 1027 1618 1030
rect 1610 1023 1614 1027
rect 1610 1017 1618 1023
rect 1623 1028 1636 1029
rect 1623 1024 1626 1028
rect 1630 1025 1636 1028
rect 1640 1028 1661 1029
rect 1640 1025 1649 1028
rect 1630 1024 1631 1025
rect 1648 1024 1649 1025
rect 1653 1025 1661 1028
rect 1674 1028 1698 1030
rect 1728 1029 1732 1030
rect 1674 1027 1694 1028
rect 1653 1024 1654 1025
rect 1623 1017 1629 1024
rect 1678 1024 1694 1027
rect 1743 1027 1749 1034
rect 1718 1026 1719 1027
rect 1678 1023 1698 1024
rect 1640 1021 1644 1022
rect 1674 1021 1698 1023
rect 1711 1023 1719 1026
rect 1723 1026 1724 1027
rect 1741 1026 1742 1027
rect 1723 1023 1742 1026
rect 1746 1023 1749 1027
rect 1711 1022 1749 1023
rect 1754 1028 1762 1034
rect 1758 1024 1762 1028
rect 1610 1013 1614 1017
rect 1640 1013 1644 1017
rect 1649 1018 1698 1021
rect 1653 1017 1698 1018
rect 1732 1019 1735 1022
rect 1649 1013 1653 1014
rect 1610 949 1618 1013
rect 1623 1009 1644 1013
rect 1656 1011 1669 1014
rect 1623 999 1627 1009
rect 1640 1008 1653 1009
rect 1656 1008 1664 1011
rect 1623 994 1627 995
rect 1631 1002 1636 1006
rect 1640 1004 1649 1008
rect 1640 1003 1653 1004
rect 1663 1007 1664 1008
rect 1668 1007 1669 1011
rect 1663 1005 1669 1007
rect 1631 998 1632 1002
rect 1663 1001 1664 1005
rect 1668 1001 1669 1005
rect 1674 1013 1698 1017
rect 1678 1009 1698 1013
rect 1732 1016 1747 1019
rect 1719 1012 1723 1013
rect 1674 999 1698 1009
rect 1631 997 1636 998
rect 1631 993 1638 997
rect 1642 993 1645 997
rect 1652 994 1653 998
rect 1657 995 1674 998
rect 1678 995 1698 999
rect 1657 994 1698 995
rect 1674 991 1698 994
rect 1674 987 1694 991
rect 1628 980 1664 983
rect 1674 975 1698 987
rect 1703 1011 1707 1012
rect 1703 989 1707 1007
rect 1711 1008 1748 1012
rect 1711 1001 1715 1008
rect 1726 1003 1727 1004
rect 1711 996 1715 997
rect 1719 1000 1727 1003
rect 1731 1003 1732 1004
rect 1731 1000 1740 1003
rect 1719 999 1740 1000
rect 1719 992 1723 999
rect 1718 991 1723 992
rect 1703 985 1712 989
rect 1722 987 1723 991
rect 1718 986 1723 987
rect 1727 994 1731 995
rect 1708 982 1712 985
rect 1727 982 1731 990
rect 1708 978 1731 982
rect 1736 983 1740 999
rect 1744 993 1748 1008
rect 1744 988 1748 989
rect 1754 1011 1762 1024
rect 1758 1007 1762 1011
rect 1736 979 1742 983
rect 1746 979 1747 983
rect 1674 971 1697 975
rect 1701 971 1704 975
rect 1708 971 1709 975
rect 1642 956 1659 959
rect 1656 951 1659 956
rect 1655 950 1669 951
rect 1610 945 1614 949
rect 1630 946 1631 950
rect 1635 946 1651 950
rect 1655 946 1656 950
rect 1660 946 1669 950
rect 1540 918 1548 940
rect 1554 935 1558 936
rect 1554 920 1558 931
rect 1561 928 1564 941
rect 1610 940 1618 945
rect 1604 937 1618 940
rect 1604 936 1627 937
rect 1573 932 1583 936
rect 1592 935 1623 936
rect 1596 934 1623 935
rect 1596 931 1604 934
rect 1592 930 1604 931
rect 1608 932 1623 934
rect 1608 931 1627 932
rect 1631 936 1637 943
rect 1647 942 1651 946
rect 1647 938 1650 942
rect 1654 938 1656 942
rect 1663 939 1669 946
rect 1631 934 1644 936
rect 1608 930 1618 931
rect 1631 930 1635 934
rect 1639 930 1644 934
rect 1561 924 1574 928
rect 1570 922 1574 924
rect 1578 923 1582 928
rect 1540 917 1551 918
rect 1540 913 1547 917
rect 1554 916 1566 920
rect 1540 912 1551 913
rect 1540 906 1548 912
rect 1540 902 1544 906
rect 1540 896 1548 902
rect 1554 905 1558 913
rect 1562 912 1566 916
rect 1585 921 1592 925
rect 1596 921 1597 925
rect 1570 915 1574 918
rect 1585 912 1589 921
rect 1604 916 1618 930
rect 1652 925 1656 938
rect 1674 932 1698 971
rect 1716 965 1720 978
rect 1728 969 1733 973
rect 1737 969 1741 973
rect 1754 972 1762 1007
rect 1799 1040 1803 1090
rect 1799 987 1804 1040
rect 1799 986 1813 987
rect 1799 982 1808 986
rect 1812 982 1813 986
rect 1728 967 1741 969
rect 1703 961 1709 964
rect 1716 961 1718 965
rect 1722 961 1725 965
rect 1703 957 1704 961
rect 1708 957 1709 961
rect 1721 957 1725 961
rect 1735 960 1741 967
rect 1745 971 1762 972
rect 1749 967 1762 971
rect 1745 966 1762 967
rect 1754 958 1762 966
rect 1703 953 1712 957
rect 1716 953 1717 957
rect 1721 953 1737 957
rect 1741 953 1742 957
rect 1758 954 1762 958
rect 1703 952 1717 953
rect 1707 938 1746 941
rect 1750 938 1751 941
rect 1663 928 1664 932
rect 1668 928 1671 932
rect 1675 928 1698 932
rect 1625 920 1626 924
rect 1630 920 1636 924
rect 1562 908 1577 912
rect 1581 908 1589 912
rect 1592 915 1618 916
rect 1596 911 1618 915
rect 1592 910 1618 911
rect 1604 906 1618 910
rect 1554 901 1556 905
rect 1560 904 1561 905
rect 1591 904 1592 905
rect 1560 901 1592 904
rect 1596 901 1599 905
rect 1554 900 1599 901
rect 1608 902 1618 906
rect 1144 894 1409 895
rect 1043 891 1451 894
rect 1059 872 1062 891
rect 1142 872 1145 891
rect 1155 883 1185 886
rect 1104 857 1108 868
rect 1087 853 1090 856
rect 1104 847 1107 857
rect 1159 852 1162 855
rect 1104 843 1105 847
rect 1176 846 1179 868
rect 1182 856 1185 883
rect 1205 872 1208 891
rect 1215 886 1218 891
rect 1259 872 1262 891
rect 1269 886 1272 891
rect 1315 872 1318 891
rect 1325 886 1328 891
rect 1369 872 1372 891
rect 1379 886 1382 891
rect 1189 863 1192 868
rect 1222 863 1225 868
rect 1189 860 1225 863
rect 1182 853 1187 856
rect 1191 852 1193 855
rect 1213 852 1214 855
rect 1222 851 1225 860
rect 1243 863 1246 868
rect 1276 863 1279 868
rect 1243 860 1279 863
rect 1299 863 1302 868
rect 1332 863 1335 868
rect 1299 860 1335 863
rect 1353 863 1356 868
rect 1386 863 1389 868
rect 1353 860 1389 863
rect 1229 851 1232 860
rect 1243 855 1250 856
rect 1243 853 1247 855
rect 1264 851 1268 854
rect 1222 848 1232 851
rect 1104 835 1107 843
rect 1176 842 1177 846
rect 1176 834 1179 842
rect 1222 835 1225 848
rect 1264 847 1267 851
rect 1276 848 1279 860
rect 1332 859 1335 860
rect 1300 852 1303 855
rect 1276 845 1295 848
rect 1276 835 1279 845
rect 1324 849 1327 851
rect 1312 841 1315 847
rect 1326 845 1327 849
rect 1324 844 1327 845
rect 1289 838 1315 841
rect 1332 835 1335 855
rect 1356 851 1357 854
rect 1375 855 1381 856
rect 1375 853 1378 855
rect 1356 842 1359 851
rect 1386 850 1389 860
rect 1358 838 1359 842
rect 1386 835 1389 846
rect 1070 825 1073 831
rect 1142 825 1145 830
rect 1188 825 1191 831
rect 1242 825 1245 831
rect 1298 825 1301 831
rect 1352 825 1355 831
rect 1002 821 1024 824
rect 700 817 868 820
rect 700 816 824 817
rect 829 813 832 817
rect 373 802 409 806
rect 413 802 423 806
rect 427 802 437 806
rect 441 803 520 806
rect 441 802 504 803
rect 189 791 211 795
rect 215 791 216 795
rect 240 794 252 795
rect 228 791 245 794
rect 189 790 193 791
rect 175 789 179 790
rect 156 786 161 789
rect 156 785 157 786
rect 86 775 89 779
rect 93 775 94 779
rect 98 775 99 779
rect 103 775 104 779
rect 109 778 113 779
rect 148 782 157 785
rect 182 786 193 790
rect 182 782 186 786
rect 200 783 201 787
rect 205 783 216 787
rect 78 774 83 775
rect 78 766 82 774
rect 98 770 104 775
rect 85 766 86 770
rect 90 766 104 770
rect 110 768 114 771
rect 148 768 151 782
rect 156 781 161 782
rect 165 780 186 782
rect 78 757 82 762
rect 78 756 83 757
rect 78 752 79 756
rect 83 752 90 755
rect 78 749 90 752
rect 94 753 98 766
rect 157 776 165 777
rect 169 778 186 780
rect 157 773 169 776
rect 110 762 114 764
rect 101 758 105 762
rect 109 758 114 762
rect 101 757 114 758
rect 157 761 161 773
rect 182 771 186 778
rect 190 776 191 780
rect 195 779 196 780
rect 195 776 207 779
rect 190 775 207 776
rect 203 772 207 775
rect 203 771 208 772
rect 171 765 177 770
rect 182 767 194 771
rect 198 767 199 771
rect 203 767 204 771
rect 171 763 173 765
rect 164 761 173 763
rect 203 766 208 767
rect 212 767 216 783
rect 203 762 207 766
rect 164 757 177 761
rect 183 758 207 762
rect 212 763 214 767
rect 157 756 161 757
rect 183 756 187 758
rect 94 749 108 753
rect 112 749 113 753
rect 170 749 171 753
rect 175 749 176 753
rect 212 754 216 763
rect 183 751 187 752
rect 192 750 193 754
rect 197 750 216 754
rect 228 751 231 791
rect 240 790 245 791
rect 249 790 252 794
rect 240 789 252 790
rect 259 794 263 797
rect 273 791 295 795
rect 299 791 300 795
rect 273 790 277 791
rect 259 789 263 790
rect 240 786 245 789
rect 240 782 241 786
rect 266 786 277 790
rect 266 782 270 786
rect 284 783 285 787
rect 289 783 300 787
rect 240 781 245 782
rect 249 780 270 782
rect 241 776 249 777
rect 253 778 270 780
rect 241 773 253 776
rect 241 761 245 773
rect 266 771 270 778
rect 274 776 275 780
rect 279 779 280 780
rect 279 776 291 779
rect 274 775 291 776
rect 287 772 291 775
rect 296 775 300 783
rect 310 780 314 787
rect 310 779 315 780
rect 310 775 311 779
rect 318 779 322 800
rect 325 794 338 795
rect 325 790 328 794
rect 332 790 334 794
rect 325 789 338 790
rect 325 782 331 789
rect 341 783 345 800
rect 355 782 370 785
rect 318 775 321 779
rect 325 775 326 779
rect 330 775 331 779
rect 335 775 336 779
rect 341 778 345 779
rect 287 771 292 772
rect 255 765 261 770
rect 266 767 278 771
rect 282 767 283 771
rect 287 767 288 771
rect 255 763 257 765
rect 248 761 257 763
rect 287 766 292 767
rect 296 771 303 775
rect 310 774 315 775
rect 287 762 291 766
rect 248 757 261 761
rect 267 758 291 762
rect 241 756 245 757
rect 267 756 271 758
rect 170 744 176 749
rect 254 749 255 753
rect 259 749 260 753
rect 296 754 300 771
rect 310 766 314 774
rect 330 770 336 775
rect 317 766 318 770
rect 322 766 336 770
rect 342 769 346 771
rect 267 751 271 752
rect 276 750 277 754
rect 281 750 300 754
rect 304 763 314 766
rect 304 751 307 763
rect 254 744 260 749
rect 310 757 314 763
rect 310 756 315 757
rect 310 752 311 756
rect 315 752 322 755
rect 310 749 322 752
rect 326 753 330 766
rect 342 762 346 765
rect 333 758 337 762
rect 341 758 346 762
rect 333 757 346 758
rect 326 749 340 753
rect 344 749 345 753
rect 77 740 80 744
rect 84 740 90 744
rect 94 740 158 744
rect 162 740 211 744
rect 215 740 242 744
rect 246 740 295 744
rect 299 740 312 744
rect 316 740 322 744
rect 326 740 345 744
rect 77 737 345 740
rect 77 736 350 737
rect 167 734 211 736
rect 167 730 173 734
rect 177 730 201 734
rect 205 730 211 734
rect 367 732 370 782
rect 171 722 177 730
rect 171 718 172 722
rect 176 718 177 722
rect 182 722 186 723
rect 191 722 197 730
rect 298 727 339 730
rect 368 728 370 732
rect 191 718 192 722
rect 196 718 197 722
rect 202 722 207 725
rect 206 718 207 722
rect 182 715 186 718
rect 202 717 207 718
rect 182 711 199 715
rect 171 699 175 709
rect 179 704 184 708
rect 195 707 199 711
rect 179 696 185 700
rect 189 696 192 700
rect 43 671 48 689
rect 179 690 183 696
rect 195 692 199 703
rect 166 687 183 690
rect 187 688 199 692
rect 203 706 207 717
rect 295 709 318 712
rect 323 709 324 712
rect 203 703 230 706
rect 187 684 191 688
rect 203 687 207 703
rect 202 686 207 687
rect 171 680 172 684
rect 176 680 191 684
rect 194 682 202 684
rect 206 682 207 686
rect 194 680 207 682
rect 224 693 230 703
rect 189 674 190 677
rect 6 669 48 671
rect 167 673 190 674
rect 194 674 195 677
rect 194 673 201 674
rect 167 670 201 673
rect 205 670 211 674
rect 167 669 211 670
rect 6 666 211 669
rect 6 665 167 666
rect 6 664 47 665
rect 6 660 12 664
rect 7 450 12 660
rect 224 597 231 693
rect 336 626 339 727
rect 348 708 364 712
rect 373 691 377 802
rect 407 782 411 789
rect 407 781 412 782
rect 407 777 408 781
rect 415 781 419 802
rect 422 796 435 797
rect 422 792 425 796
rect 429 792 431 796
rect 422 791 435 792
rect 422 784 428 791
rect 438 785 442 802
rect 508 802 520 803
rect 524 803 604 806
rect 524 802 588 803
rect 485 791 497 797
rect 504 796 508 799
rect 592 802 604 803
rect 608 802 641 806
rect 645 802 655 806
rect 659 802 669 806
rect 673 802 679 806
rect 693 806 697 809
rect 700 809 1006 813
rect 518 793 540 797
rect 544 793 545 797
rect 569 796 581 797
rect 518 792 522 793
rect 504 791 508 792
rect 485 788 490 791
rect 485 787 486 788
rect 415 777 418 781
rect 422 777 423 781
rect 427 777 428 781
rect 432 777 433 781
rect 438 780 442 781
rect 477 784 486 787
rect 511 788 522 792
rect 569 792 574 796
rect 578 792 581 796
rect 569 791 581 792
rect 588 796 592 799
rect 602 793 624 797
rect 628 793 629 797
rect 602 792 606 793
rect 588 791 592 792
rect 511 784 515 788
rect 529 785 530 789
rect 534 785 545 789
rect 407 776 412 777
rect 407 768 411 776
rect 427 772 433 777
rect 414 768 415 772
rect 419 768 433 772
rect 439 770 443 773
rect 407 759 411 764
rect 407 758 412 759
rect 407 754 408 758
rect 412 754 419 757
rect 407 751 419 754
rect 423 755 427 768
rect 439 764 443 766
rect 430 760 434 764
rect 438 760 443 764
rect 430 759 443 760
rect 423 751 437 755
rect 441 751 442 755
rect 467 753 470 773
rect 477 770 480 784
rect 485 783 490 784
rect 494 782 515 784
rect 486 778 494 779
rect 498 780 515 782
rect 486 775 498 778
rect 486 763 490 775
rect 511 773 515 780
rect 519 778 520 782
rect 524 781 525 782
rect 524 778 536 781
rect 519 777 536 778
rect 532 774 536 777
rect 532 773 537 774
rect 500 767 506 772
rect 511 769 523 773
rect 527 769 528 773
rect 532 769 533 773
rect 500 765 502 767
rect 493 763 502 765
rect 532 768 537 769
rect 541 769 545 785
rect 569 788 574 791
rect 569 784 570 788
rect 595 788 606 792
rect 595 784 599 788
rect 613 785 614 789
rect 618 785 629 789
rect 569 783 574 784
rect 578 782 599 784
rect 570 778 578 779
rect 582 780 599 782
rect 570 775 582 778
rect 532 764 536 768
rect 493 759 506 763
rect 512 760 536 764
rect 541 765 543 769
rect 486 758 490 759
rect 512 758 516 760
rect 499 751 500 755
rect 504 751 505 755
rect 541 756 545 765
rect 570 763 574 775
rect 595 773 599 780
rect 603 778 604 782
rect 608 781 609 782
rect 608 778 620 781
rect 603 777 620 778
rect 616 774 620 777
rect 625 780 629 785
rect 639 782 643 789
rect 639 781 644 782
rect 625 777 632 780
rect 639 777 640 781
rect 647 781 651 802
rect 654 796 667 797
rect 654 792 657 796
rect 661 792 663 796
rect 654 791 667 792
rect 654 784 660 791
rect 670 785 674 802
rect 647 777 650 781
rect 654 777 655 781
rect 659 777 660 781
rect 664 777 665 781
rect 670 780 674 781
rect 616 773 621 774
rect 584 767 590 772
rect 595 769 607 773
rect 611 769 612 773
rect 616 769 617 773
rect 584 765 586 767
rect 577 763 586 765
rect 616 768 621 769
rect 616 764 620 768
rect 577 759 590 763
rect 596 760 620 764
rect 570 758 574 759
rect 596 758 600 760
rect 512 753 516 754
rect 521 752 522 756
rect 526 752 545 756
rect 499 746 505 751
rect 583 751 584 755
rect 588 751 589 755
rect 625 756 629 777
rect 639 776 644 777
rect 639 768 643 776
rect 659 772 665 777
rect 646 768 647 772
rect 651 768 665 772
rect 671 771 675 773
rect 596 753 600 754
rect 605 752 606 756
rect 610 752 629 756
rect 633 765 643 768
rect 633 753 636 765
rect 583 746 589 751
rect 639 759 643 765
rect 639 758 644 759
rect 639 754 640 758
rect 644 754 651 757
rect 639 751 651 754
rect 655 755 659 768
rect 693 770 696 806
rect 671 764 675 767
rect 662 760 666 764
rect 670 760 675 764
rect 662 759 675 760
rect 691 763 696 770
rect 700 805 736 809
rect 740 805 750 809
rect 754 805 764 809
rect 768 806 847 809
rect 768 805 831 806
rect 655 751 669 755
rect 673 751 674 755
rect 406 742 409 746
rect 413 742 419 746
rect 423 742 487 746
rect 491 742 540 746
rect 544 742 571 746
rect 575 742 624 746
rect 628 742 641 746
rect 645 742 651 746
rect 655 742 679 746
rect 387 739 672 742
rect 406 738 672 739
rect 676 738 679 742
rect 496 736 540 738
rect 496 732 502 736
rect 506 732 530 736
rect 534 732 540 736
rect 395 728 416 731
rect 372 671 377 691
rect 412 693 415 728
rect 467 727 470 729
rect 500 724 506 732
rect 467 709 470 723
rect 500 720 501 724
rect 505 720 506 724
rect 511 724 515 725
rect 520 724 526 732
rect 666 727 670 728
rect 691 727 695 763
rect 520 720 521 724
rect 525 720 526 724
rect 531 724 536 727
rect 535 720 536 724
rect 666 724 695 727
rect 666 723 693 724
rect 511 717 515 720
rect 531 719 536 720
rect 511 713 528 717
rect 439 705 467 708
rect 412 690 432 693
rect 429 681 432 690
rect 426 679 432 681
rect 430 677 432 679
rect 439 679 443 705
rect 500 701 504 711
rect 508 706 513 710
rect 524 709 528 713
rect 508 698 514 702
rect 518 698 521 702
rect 508 692 512 698
rect 524 694 528 705
rect 495 689 512 692
rect 516 690 528 694
rect 516 686 520 690
rect 532 689 536 719
rect 563 715 645 720
rect 666 700 670 723
rect 531 688 536 689
rect 500 682 501 686
rect 505 682 520 686
rect 523 684 531 686
rect 535 686 536 688
rect 535 684 540 686
rect 523 682 540 684
rect 518 676 519 679
rect 496 675 519 676
rect 523 676 524 679
rect 523 675 530 676
rect 496 672 530 675
rect 534 672 540 676
rect 496 671 540 672
rect 372 668 540 671
rect 372 667 420 668
rect 438 667 444 668
rect 462 667 496 668
rect 432 661 450 664
rect 485 660 489 667
rect 368 658 412 660
rect 461 658 505 660
rect 548 658 592 660
rect 368 656 592 658
rect 368 652 374 656
rect 378 655 467 656
rect 378 652 412 655
rect 461 652 467 655
rect 471 655 554 656
rect 471 652 505 655
rect 548 652 554 655
rect 558 652 592 656
rect 382 644 388 652
rect 382 640 383 644
rect 387 640 388 644
rect 393 646 397 647
rect 402 646 408 652
rect 443 646 454 649
rect 402 642 403 646
rect 407 642 408 646
rect 372 639 377 640
rect 372 635 373 639
rect 393 639 397 642
rect 372 632 377 635
rect 372 628 373 632
rect 372 627 377 628
rect 380 635 393 637
rect 380 633 397 635
rect 404 635 435 639
rect 372 626 376 627
rect 336 622 376 626
rect 372 609 376 622
rect 380 622 384 633
rect 395 626 400 630
rect 404 626 408 635
rect 387 618 390 622
rect 394 618 401 622
rect 380 614 384 618
rect 380 610 392 614
rect 396 613 401 618
rect 372 608 377 609
rect 372 604 373 608
rect 377 604 384 607
rect 372 601 384 604
rect 388 606 392 610
rect 395 609 411 613
rect 388 602 403 606
rect 407 602 408 606
rect 431 602 435 635
rect 451 636 454 646
rect 475 644 481 652
rect 475 640 476 644
rect 480 640 481 644
rect 486 646 490 647
rect 495 646 501 652
rect 495 642 496 646
rect 500 642 501 646
rect 562 644 568 652
rect 541 643 557 644
rect 465 639 470 640
rect 465 636 466 639
rect 451 635 466 636
rect 486 639 490 642
rect 451 633 470 635
rect 465 632 470 633
rect 465 628 466 632
rect 465 627 470 628
rect 473 635 486 637
rect 473 633 490 635
rect 465 609 469 627
rect 473 622 477 633
rect 497 630 501 639
rect 545 639 557 643
rect 562 640 563 644
rect 567 640 568 644
rect 573 646 577 647
rect 582 646 588 652
rect 582 642 583 646
rect 587 642 588 646
rect 545 638 553 639
rect 552 635 553 638
rect 573 639 577 642
rect 552 632 557 635
rect 488 626 493 630
rect 497 626 508 630
rect 552 628 553 632
rect 552 627 557 628
rect 560 635 573 637
rect 560 633 577 635
rect 480 618 483 622
rect 487 618 494 622
rect 473 614 477 618
rect 473 610 485 614
rect 465 608 470 609
rect 465 604 466 608
rect 470 604 477 607
rect 465 601 477 604
rect 481 606 485 610
rect 489 613 494 618
rect 489 609 504 613
rect 552 609 556 627
rect 560 622 564 633
rect 584 630 588 639
rect 575 626 580 630
rect 584 626 597 630
rect 628 622 632 660
rect 665 662 670 700
rect 700 694 704 805
rect 734 785 738 792
rect 734 784 739 785
rect 734 780 735 784
rect 742 784 746 805
rect 749 799 762 800
rect 749 795 752 799
rect 756 795 758 799
rect 749 794 762 795
rect 749 787 755 794
rect 765 788 769 805
rect 835 805 847 806
rect 851 806 931 809
rect 851 805 915 806
rect 812 794 824 800
rect 831 799 835 802
rect 919 805 931 806
rect 935 805 968 809
rect 972 805 982 809
rect 986 805 996 809
rect 1000 805 1006 809
rect 845 796 867 800
rect 871 796 872 800
rect 896 799 908 800
rect 845 795 849 796
rect 831 794 835 795
rect 812 791 817 794
rect 812 790 813 791
rect 742 780 745 784
rect 749 780 750 784
rect 754 780 755 784
rect 759 780 760 784
rect 765 783 769 784
rect 804 787 813 790
rect 838 791 849 795
rect 896 795 901 799
rect 905 795 908 799
rect 896 794 908 795
rect 915 799 919 802
rect 929 796 951 800
rect 955 796 956 800
rect 929 795 933 796
rect 915 794 919 795
rect 838 787 842 791
rect 856 788 857 792
rect 861 788 872 792
rect 734 779 739 780
rect 734 771 738 779
rect 754 775 760 780
rect 741 771 742 775
rect 746 771 760 775
rect 766 773 770 776
rect 804 773 807 787
rect 812 786 817 787
rect 821 785 842 787
rect 734 762 738 767
rect 734 761 739 762
rect 734 757 735 761
rect 739 757 746 760
rect 734 754 746 757
rect 750 758 754 771
rect 813 781 821 782
rect 825 783 842 785
rect 813 778 825 781
rect 766 767 770 769
rect 757 763 761 767
rect 765 763 770 767
rect 757 762 770 763
rect 813 766 817 778
rect 838 776 842 783
rect 846 781 847 785
rect 851 784 852 785
rect 851 781 863 784
rect 846 780 863 781
rect 859 777 863 780
rect 859 776 864 777
rect 827 770 833 775
rect 838 772 850 776
rect 854 772 855 776
rect 859 772 860 776
rect 827 768 829 770
rect 813 761 817 762
rect 820 766 829 768
rect 859 771 864 772
rect 868 772 872 788
rect 896 791 901 794
rect 896 787 897 791
rect 922 791 933 795
rect 922 787 926 791
rect 940 788 941 792
rect 945 788 956 792
rect 896 786 901 787
rect 905 785 926 787
rect 897 781 905 782
rect 909 783 926 785
rect 897 778 909 781
rect 859 767 863 771
rect 820 762 833 766
rect 839 763 863 767
rect 868 768 870 772
rect 750 754 764 758
rect 768 754 769 758
rect 820 757 823 762
rect 839 761 843 763
rect 809 753 823 757
rect 826 754 827 758
rect 831 754 832 758
rect 868 759 872 768
rect 897 766 901 778
rect 922 776 926 783
rect 930 781 931 785
rect 935 784 936 785
rect 935 781 947 784
rect 930 780 947 781
rect 943 777 947 780
rect 952 782 956 788
rect 966 785 970 792
rect 966 784 971 785
rect 952 779 959 782
rect 966 780 967 784
rect 974 784 978 805
rect 981 799 994 800
rect 981 795 984 799
rect 988 795 990 799
rect 981 794 994 795
rect 981 787 987 794
rect 997 788 1001 805
rect 974 780 977 784
rect 981 780 982 784
rect 986 780 987 784
rect 991 780 992 784
rect 997 783 1001 784
rect 966 779 971 780
rect 943 776 948 777
rect 911 770 917 775
rect 922 772 934 776
rect 938 772 939 776
rect 943 772 944 776
rect 911 768 913 770
rect 904 766 913 768
rect 943 771 948 772
rect 943 767 947 771
rect 904 762 917 766
rect 923 763 947 767
rect 897 761 901 762
rect 923 761 927 763
rect 839 756 843 757
rect 848 755 849 759
rect 853 755 872 759
rect 809 749 813 753
rect 826 749 832 754
rect 910 754 911 758
rect 915 754 916 758
rect 952 759 956 779
rect 966 771 970 779
rect 986 775 992 780
rect 973 771 974 775
rect 978 771 992 775
rect 998 774 1002 776
rect 923 756 927 757
rect 932 755 933 759
rect 937 755 956 759
rect 960 768 970 771
rect 960 756 963 768
rect 910 749 916 754
rect 966 762 970 768
rect 966 761 971 762
rect 966 757 967 761
rect 971 757 978 760
rect 966 754 978 757
rect 982 758 986 771
rect 998 767 1002 770
rect 989 763 993 767
rect 997 763 1002 767
rect 989 762 1002 763
rect 982 754 996 758
rect 1000 754 1001 758
rect 733 746 736 749
rect 732 745 736 746
rect 740 745 746 749
rect 750 745 814 749
rect 818 745 867 749
rect 871 745 898 749
rect 902 745 951 749
rect 955 745 968 749
rect 972 745 978 749
rect 982 745 1006 749
rect 732 743 1006 745
rect 713 742 1006 743
rect 716 741 1006 742
rect 716 740 735 741
rect 823 739 867 741
rect 823 735 829 739
rect 833 735 857 739
rect 861 735 867 739
rect 770 733 774 734
rect 714 715 743 720
rect 699 674 704 694
rect 770 692 774 729
rect 827 727 833 735
rect 827 723 828 727
rect 832 723 833 727
rect 838 727 842 728
rect 847 727 853 735
rect 847 723 848 727
rect 852 723 853 727
rect 858 727 863 730
rect 862 723 863 727
rect 838 720 842 723
rect 858 722 863 723
rect 838 716 855 720
rect 827 704 831 714
rect 835 709 840 713
rect 851 712 855 716
rect 835 701 841 705
rect 845 701 848 705
rect 835 695 839 701
rect 851 697 855 708
rect 822 692 839 695
rect 843 693 855 697
rect 859 717 875 722
rect 843 689 847 693
rect 859 692 863 717
rect 858 691 863 692
rect 827 685 828 689
rect 832 685 847 689
rect 850 687 858 689
rect 862 687 863 691
rect 850 685 863 687
rect 845 679 846 682
rect 823 678 846 679
rect 850 679 851 682
rect 850 678 857 679
rect 823 675 857 678
rect 861 675 867 679
rect 823 674 867 675
rect 699 671 867 674
rect 699 670 823 671
rect 1021 666 1024 821
rect 1030 822 1391 825
rect 1030 683 1033 822
rect 1214 819 1219 822
rect 1320 819 1324 822
rect 1146 816 1395 819
rect 1146 811 1149 816
rect 1192 810 1195 816
rect 1246 810 1249 816
rect 1302 810 1305 816
rect 1356 810 1359 816
rect 1180 799 1183 807
rect 1180 795 1181 799
rect 1163 786 1166 789
rect 1180 773 1183 795
rect 1226 793 1229 806
rect 1226 790 1236 793
rect 1268 790 1271 794
rect 1280 796 1283 806
rect 1280 793 1299 796
rect 1328 796 1331 797
rect 1195 786 1197 789
rect 1217 786 1218 789
rect 1226 781 1229 790
rect 1193 778 1229 781
rect 1193 773 1196 778
rect 1226 773 1229 778
rect 1233 781 1236 790
rect 1247 786 1251 788
rect 1268 787 1272 790
rect 1247 785 1254 786
rect 1280 781 1283 793
rect 1330 792 1331 796
rect 1328 790 1331 792
rect 1304 786 1307 789
rect 1336 786 1339 806
rect 1362 799 1363 803
rect 1360 790 1363 799
rect 1390 795 1393 806
rect 1360 787 1361 790
rect 1379 786 1382 788
rect 1379 785 1385 786
rect 1336 781 1339 782
rect 1390 781 1393 791
rect 1247 778 1283 781
rect 1247 773 1250 778
rect 1280 773 1283 778
rect 1303 778 1339 781
rect 1303 773 1306 778
rect 1336 773 1339 778
rect 1357 778 1393 781
rect 1357 773 1360 778
rect 1390 773 1393 778
rect 1146 752 1149 769
rect 1209 752 1212 769
rect 1219 752 1222 755
rect 1263 752 1266 769
rect 1273 752 1276 755
rect 1319 752 1322 769
rect 1329 752 1332 755
rect 1373 752 1376 769
rect 1404 759 1409 891
rect 1415 890 1462 891
rect 1415 886 1421 890
rect 1425 886 1431 890
rect 1435 886 1462 890
rect 1434 880 1447 881
rect 1434 876 1442 880
rect 1446 876 1447 880
rect 1442 873 1447 876
rect 1419 868 1420 872
rect 1424 868 1439 872
rect 1446 869 1447 873
rect 1442 868 1447 869
rect 1417 861 1423 865
rect 1419 857 1423 861
rect 1419 856 1431 857
rect 1419 852 1423 856
rect 1427 852 1431 856
rect 1419 851 1431 852
rect 1435 856 1439 868
rect 1435 847 1439 852
rect 1443 855 1447 868
rect 1541 880 1547 896
rect 1563 895 1566 900
rect 1604 896 1618 902
rect 1610 892 1614 896
rect 1541 874 1557 880
rect 1610 879 1618 892
rect 1624 914 1628 915
rect 1624 895 1628 910
rect 1632 904 1636 920
rect 1641 921 1664 925
rect 1641 913 1645 921
rect 1660 918 1664 921
rect 1641 908 1645 909
rect 1649 916 1654 917
rect 1649 912 1650 916
rect 1660 914 1669 918
rect 1649 911 1654 912
rect 1649 904 1653 911
rect 1632 903 1653 904
rect 1632 900 1641 903
rect 1640 899 1641 900
rect 1645 900 1653 903
rect 1657 906 1661 907
rect 1645 899 1646 900
rect 1657 895 1661 902
rect 1624 893 1661 895
rect 1624 891 1637 893
rect 1641 891 1661 893
rect 1665 896 1669 914
rect 1665 891 1669 892
rect 1674 916 1698 928
rect 1678 912 1698 916
rect 1674 907 1698 912
rect 1674 903 1694 907
rect 1674 891 1698 903
rect 1703 927 1707 928
rect 1703 905 1707 923
rect 1711 926 1731 928
rect 1735 926 1748 928
rect 1711 924 1748 926
rect 1711 917 1715 924
rect 1726 919 1727 920
rect 1711 912 1715 913
rect 1719 916 1727 919
rect 1731 919 1732 920
rect 1731 916 1740 919
rect 1719 915 1740 916
rect 1719 908 1723 915
rect 1718 907 1723 908
rect 1703 901 1712 905
rect 1722 903 1723 907
rect 1718 902 1723 903
rect 1727 910 1731 911
rect 1708 898 1712 901
rect 1727 898 1731 906
rect 1708 894 1731 898
rect 1736 899 1740 915
rect 1744 909 1748 924
rect 1744 904 1748 905
rect 1754 927 1762 954
rect 1772 938 1788 941
rect 1758 923 1762 927
rect 1754 917 1768 923
rect 1785 919 1788 938
rect 1754 913 1764 917
rect 1773 918 1818 919
rect 1773 914 1776 918
rect 1780 915 1812 918
rect 1780 914 1781 915
rect 1811 914 1812 915
rect 1816 914 1818 918
rect 1754 909 1768 913
rect 1754 908 1780 909
rect 1754 904 1776 908
rect 1754 903 1780 904
rect 1783 907 1791 911
rect 1795 907 1810 911
rect 1736 895 1742 899
rect 1746 895 1747 899
rect 1576 875 1618 879
rect 1443 852 1492 855
rect 1443 848 1447 852
rect 1419 843 1420 847
rect 1424 843 1439 847
rect 1442 847 1447 848
rect 1446 843 1447 847
rect 1442 840 1447 843
rect 1430 835 1431 839
rect 1435 835 1436 839
rect 1446 836 1447 840
rect 1442 835 1447 836
rect 1430 830 1436 835
rect 1415 827 1421 830
rect 1416 826 1421 827
rect 1425 826 1457 830
rect 1416 824 1457 826
rect 1416 823 1469 824
rect 1415 822 1469 823
rect 1416 821 1469 822
rect 1416 817 1422 821
rect 1426 820 1469 821
rect 1426 817 1457 820
rect 1431 812 1437 817
rect 1431 808 1432 812
rect 1436 808 1437 812
rect 1443 811 1448 812
rect 1447 807 1448 811
rect 1443 804 1448 807
rect 1420 800 1421 804
rect 1425 800 1440 804
rect 1420 795 1432 796
rect 1420 791 1424 795
rect 1428 791 1432 795
rect 1420 790 1432 791
rect 1436 795 1440 800
rect 1447 800 1448 804
rect 1443 799 1448 800
rect 1420 786 1424 790
rect 1419 782 1424 786
rect 1436 779 1440 791
rect 1444 787 1448 799
rect 1444 783 1447 787
rect 1444 779 1448 783
rect 1420 775 1421 779
rect 1425 775 1440 779
rect 1443 778 1448 779
rect 1447 774 1448 778
rect 1443 771 1448 774
rect 1435 767 1443 771
rect 1447 767 1448 771
rect 1435 766 1448 767
rect 1416 759 1422 761
rect 1404 757 1422 759
rect 1426 757 1432 761
rect 1436 757 1451 761
rect 1404 756 1451 757
rect 1383 752 1386 755
rect 1404 752 1409 756
rect 1042 749 1409 752
rect 1058 730 1061 749
rect 1141 747 1409 749
rect 1415 750 1451 756
rect 1092 742 1093 745
rect 1092 715 1095 742
rect 1103 732 1107 734
rect 1141 730 1144 747
rect 1152 738 1184 741
rect 1086 711 1089 714
rect 1093 712 1095 715
rect 1103 715 1107 726
rect 1103 705 1106 715
rect 1158 710 1161 713
rect 1103 701 1104 705
rect 1175 704 1178 726
rect 1181 714 1184 738
rect 1204 730 1207 747
rect 1214 744 1217 747
rect 1258 730 1261 747
rect 1268 744 1271 747
rect 1314 730 1317 747
rect 1324 744 1327 747
rect 1368 730 1371 747
rect 1378 744 1381 747
rect 1188 721 1191 726
rect 1221 721 1224 726
rect 1188 718 1224 721
rect 1181 711 1186 714
rect 1190 710 1192 713
rect 1212 710 1213 713
rect 1221 709 1224 718
rect 1242 721 1245 726
rect 1275 721 1278 726
rect 1242 718 1278 721
rect 1298 721 1301 726
rect 1331 721 1334 726
rect 1298 718 1334 721
rect 1352 721 1355 726
rect 1385 721 1388 726
rect 1352 718 1388 721
rect 1228 709 1231 718
rect 1242 713 1249 714
rect 1242 711 1246 713
rect 1263 709 1267 712
rect 1221 706 1231 709
rect 1103 693 1106 701
rect 1175 700 1176 704
rect 1175 692 1178 700
rect 1221 693 1224 706
rect 1263 705 1266 709
rect 1275 706 1278 718
rect 1331 717 1334 718
rect 1299 710 1302 713
rect 1275 703 1294 706
rect 1275 693 1278 703
rect 1323 707 1326 709
rect 1311 699 1314 705
rect 1325 703 1326 707
rect 1323 702 1326 703
rect 1288 696 1314 699
rect 1331 693 1334 713
rect 1355 709 1356 712
rect 1374 713 1380 714
rect 1374 711 1377 713
rect 1355 700 1358 709
rect 1385 708 1388 718
rect 1357 696 1358 700
rect 1385 693 1388 704
rect 1069 683 1072 689
rect 1141 683 1144 688
rect 1187 683 1190 689
rect 1241 683 1244 689
rect 1297 683 1300 689
rect 1351 683 1354 689
rect 1029 680 1390 683
rect 1213 677 1218 680
rect 1319 677 1323 680
rect 1145 674 1394 677
rect 1145 669 1148 674
rect 1083 666 1087 667
rect 1021 663 1088 666
rect 1191 668 1194 674
rect 1245 668 1248 674
rect 1301 668 1304 674
rect 1355 668 1358 674
rect 665 637 669 662
rect 947 657 951 658
rect 725 653 951 657
rect 947 649 951 653
rect 947 647 1058 649
rect 1063 647 1066 649
rect 947 644 1066 647
rect 665 636 788 637
rect 665 635 1034 636
rect 665 632 1050 635
rect 1063 628 1066 644
rect 1058 625 1066 628
rect 567 618 570 622
rect 574 618 581 622
rect 628 618 1033 622
rect 560 614 564 618
rect 560 610 572 614
rect 552 608 557 609
rect 481 602 496 606
rect 500 602 501 606
rect 552 604 553 608
rect 557 604 564 607
rect 552 601 564 604
rect 568 606 572 610
rect 576 612 581 618
rect 576 609 589 612
rect 594 610 1042 613
rect 1083 611 1087 663
rect 1179 657 1182 665
rect 1179 653 1180 657
rect 1162 644 1165 647
rect 1136 632 1139 633
rect 1106 629 1139 632
rect 1179 631 1182 653
rect 1225 651 1228 664
rect 1225 648 1235 651
rect 1267 648 1270 652
rect 1279 654 1282 664
rect 1279 651 1298 654
rect 1327 654 1330 655
rect 1194 644 1196 647
rect 1216 644 1217 647
rect 1225 639 1228 648
rect 1192 636 1228 639
rect 1192 631 1195 636
rect 1225 631 1228 636
rect 1232 639 1235 648
rect 1246 644 1250 646
rect 1267 645 1271 648
rect 1246 643 1253 644
rect 1279 639 1282 651
rect 1329 650 1330 654
rect 1327 648 1330 650
rect 1303 644 1306 647
rect 1335 644 1338 664
rect 1361 657 1362 661
rect 1359 648 1362 657
rect 1389 653 1392 664
rect 1359 645 1360 648
rect 1378 644 1381 646
rect 1378 643 1384 644
rect 1335 639 1338 640
rect 1389 639 1392 649
rect 1246 636 1282 639
rect 1246 631 1249 636
rect 1279 631 1282 636
rect 1302 636 1338 639
rect 1302 631 1305 636
rect 1335 631 1338 636
rect 1356 636 1392 639
rect 1356 631 1359 636
rect 1389 631 1392 636
rect 1136 625 1139 629
rect 1101 621 1139 625
rect 1101 618 1104 621
rect 1131 613 1134 616
rect 1139 613 1140 616
rect 1131 611 1140 613
rect 1083 607 1140 611
rect 1145 608 1148 627
rect 1208 608 1211 627
rect 1218 608 1221 613
rect 1262 608 1265 627
rect 1272 608 1275 613
rect 1318 608 1321 627
rect 1328 608 1331 613
rect 1372 608 1375 627
rect 1382 608 1385 613
rect 1403 608 1408 747
rect 1415 746 1421 750
rect 1425 746 1431 750
rect 1435 746 1451 750
rect 1434 740 1447 741
rect 1434 736 1442 740
rect 1446 736 1447 740
rect 1442 733 1447 736
rect 1419 728 1420 732
rect 1424 728 1439 732
rect 1446 729 1447 733
rect 1442 728 1447 729
rect 1419 717 1423 725
rect 1419 716 1431 717
rect 1419 712 1423 716
rect 1427 712 1431 716
rect 1419 711 1431 712
rect 1435 716 1439 728
rect 1435 707 1439 712
rect 1443 720 1447 728
rect 1443 716 1446 720
rect 1443 708 1447 716
rect 1419 703 1420 707
rect 1424 703 1439 707
rect 1442 707 1447 708
rect 1446 703 1447 707
rect 1442 700 1447 703
rect 1430 695 1431 699
rect 1435 695 1436 699
rect 1446 696 1447 700
rect 1442 695 1447 696
rect 1430 690 1436 695
rect 1454 690 1457 817
rect 1415 686 1421 690
rect 1425 686 1457 690
rect 1415 682 1457 686
rect 1438 654 1442 675
rect 1480 656 1484 852
rect 568 602 583 606
rect 587 602 588 606
rect 1143 605 1408 608
rect 1422 651 1442 654
rect 1422 607 1426 651
rect 1481 646 1484 656
rect 1541 721 1547 874
rect 1576 845 1581 875
rect 1557 841 1581 845
rect 1557 792 1561 841
rect 1576 840 1581 841
rect 1610 865 1618 875
rect 1674 887 1697 891
rect 1701 887 1704 891
rect 1708 887 1709 891
rect 1655 866 1669 867
rect 1610 861 1614 865
rect 1630 862 1631 866
rect 1635 862 1651 866
rect 1655 862 1656 866
rect 1660 862 1669 866
rect 1610 853 1618 861
rect 1610 852 1627 853
rect 1610 848 1623 852
rect 1610 847 1627 848
rect 1631 852 1637 859
rect 1647 858 1651 862
rect 1663 858 1664 862
rect 1668 858 1669 862
rect 1647 854 1650 858
rect 1654 854 1656 858
rect 1663 855 1669 858
rect 1631 850 1644 852
rect 1558 787 1561 792
rect 1584 777 1588 813
rect 1559 773 1588 777
rect 1596 733 1599 823
rect 1603 792 1606 810
rect 1610 812 1618 847
rect 1631 846 1635 850
rect 1639 846 1644 850
rect 1652 841 1656 854
rect 1674 848 1698 887
rect 1716 881 1720 894
rect 1754 889 1768 903
rect 1783 898 1787 907
rect 1798 901 1802 904
rect 1775 894 1776 898
rect 1780 894 1787 898
rect 1806 903 1810 907
rect 1814 906 1818 914
rect 1824 917 1832 923
rect 1828 913 1832 917
rect 1824 907 1832 913
rect 1821 906 1832 907
rect 1806 899 1818 903
rect 1825 902 1832 906
rect 1821 901 1832 902
rect 1790 891 1794 896
rect 1798 895 1802 897
rect 1798 891 1811 895
rect 1728 885 1733 889
rect 1737 885 1741 889
rect 1754 888 1764 889
rect 1728 883 1741 885
rect 1703 873 1709 880
rect 1716 877 1718 881
rect 1722 877 1725 881
rect 1721 873 1725 877
rect 1735 876 1741 883
rect 1745 887 1764 888
rect 1749 885 1764 887
rect 1768 888 1780 889
rect 1768 885 1776 888
rect 1749 884 1776 885
rect 1749 883 1780 884
rect 1789 883 1799 887
rect 1745 882 1768 883
rect 1754 879 1768 882
rect 1754 874 1762 879
rect 1808 878 1811 891
rect 1814 888 1818 899
rect 1814 883 1818 884
rect 1824 879 1832 901
rect 1703 869 1712 873
rect 1716 869 1717 873
rect 1721 869 1737 873
rect 1741 869 1742 873
rect 1758 870 1762 874
rect 1703 868 1717 869
rect 1713 863 1716 868
rect 1713 860 1730 863
rect 1663 844 1664 848
rect 1668 844 1671 848
rect 1675 844 1698 848
rect 1625 836 1626 840
rect 1630 836 1636 840
rect 1610 808 1614 812
rect 1610 795 1618 808
rect 1624 830 1628 831
rect 1624 811 1628 826
rect 1632 820 1636 836
rect 1641 837 1664 841
rect 1641 829 1645 837
rect 1660 834 1664 837
rect 1641 824 1645 825
rect 1649 832 1654 833
rect 1649 828 1650 832
rect 1660 830 1669 834
rect 1649 827 1654 828
rect 1649 820 1653 827
rect 1632 819 1653 820
rect 1632 816 1641 819
rect 1640 815 1641 816
rect 1645 816 1653 819
rect 1657 822 1661 823
rect 1645 815 1646 816
rect 1657 811 1661 818
rect 1624 807 1661 811
rect 1665 812 1669 830
rect 1665 807 1669 808
rect 1674 832 1698 844
rect 1678 828 1698 832
rect 1674 825 1698 828
rect 1754 853 1762 870
rect 1674 824 1715 825
rect 1674 820 1694 824
rect 1698 821 1715 824
rect 1719 821 1720 825
rect 1727 822 1730 826
rect 1734 822 1741 826
rect 1736 821 1741 822
rect 1674 810 1698 820
rect 1648 804 1651 807
rect 1625 800 1640 803
rect 1674 806 1694 810
rect 1674 802 1698 806
rect 1703 814 1704 818
rect 1708 814 1709 818
rect 1740 817 1741 821
rect 1703 812 1709 814
rect 1703 808 1704 812
rect 1708 811 1709 812
rect 1719 815 1732 816
rect 1723 811 1732 815
rect 1736 813 1741 817
rect 1745 824 1749 825
rect 1708 808 1716 811
rect 1719 810 1732 811
rect 1745 810 1749 820
rect 1703 805 1716 808
rect 1728 806 1749 810
rect 1754 806 1768 853
rect 1791 840 1818 841
rect 1791 838 1815 840
rect 1719 805 1723 806
rect 1674 801 1719 802
rect 1637 797 1640 800
rect 1674 798 1723 801
rect 1728 802 1732 806
rect 1758 802 1768 806
rect 1610 791 1614 795
rect 1610 785 1618 791
rect 1623 796 1661 797
rect 1623 792 1626 796
rect 1630 793 1649 796
rect 1630 792 1631 793
rect 1648 792 1649 793
rect 1653 793 1661 796
rect 1674 796 1698 798
rect 1728 797 1732 798
rect 1674 795 1694 796
rect 1653 792 1654 793
rect 1623 785 1629 792
rect 1678 792 1694 795
rect 1743 795 1749 802
rect 1718 794 1719 795
rect 1678 791 1698 792
rect 1640 789 1644 790
rect 1674 789 1698 791
rect 1711 791 1719 794
rect 1723 794 1724 795
rect 1741 794 1742 795
rect 1723 791 1732 794
rect 1711 790 1732 791
rect 1736 791 1742 794
rect 1746 791 1749 795
rect 1736 790 1749 791
rect 1754 796 1768 802
rect 1758 792 1768 796
rect 1754 789 1768 792
rect 1610 781 1614 785
rect 1640 781 1644 785
rect 1649 786 1698 789
rect 1653 785 1698 786
rect 1649 781 1653 782
rect 1610 757 1618 781
rect 1623 777 1644 781
rect 1656 779 1669 782
rect 1623 767 1627 777
rect 1640 776 1653 777
rect 1656 776 1664 779
rect 1623 762 1627 763
rect 1631 770 1636 774
rect 1640 772 1649 776
rect 1640 771 1653 772
rect 1663 775 1664 776
rect 1668 775 1669 779
rect 1663 773 1669 775
rect 1631 766 1632 770
rect 1663 769 1664 773
rect 1668 769 1669 773
rect 1674 781 1698 785
rect 1678 777 1698 781
rect 1674 767 1698 777
rect 1758 775 1768 789
rect 1758 772 1760 775
rect 1631 765 1636 766
rect 1631 761 1639 765
rect 1643 761 1645 765
rect 1652 762 1653 766
rect 1657 763 1674 766
rect 1678 763 1698 767
rect 1657 762 1698 763
rect 1674 760 1698 762
rect 1829 760 1833 879
rect 1674 759 1833 760
rect 1674 757 1834 759
rect 1554 732 1599 733
rect 1558 729 1599 732
rect 1612 729 1617 757
rect 1690 756 1834 757
rect 1809 755 1834 756
rect 1612 728 1738 729
rect 1612 723 1733 728
rect 1758 727 1763 732
rect 1740 722 1763 727
rect 1735 721 1763 722
rect 1541 703 1545 721
rect 1758 720 1763 721
rect 1758 717 1762 720
rect 1569 712 1590 716
rect 1552 703 1565 704
rect 1541 702 1694 703
rect 1758 702 1763 717
rect 1769 705 1772 741
rect 1541 699 1700 702
rect 1435 643 1485 646
rect 225 591 231 597
rect 230 584 231 591
rect 368 592 374 596
rect 378 592 384 596
rect 388 592 412 596
rect 461 592 467 596
rect 471 592 477 596
rect 481 592 505 596
rect 362 591 505 592
rect 548 592 554 596
rect 558 592 564 596
rect 568 592 592 596
rect 548 591 592 592
rect 362 589 592 591
rect 368 588 412 589
rect 461 588 592 589
rect 1024 589 1091 592
rect 1435 591 1439 643
rect 1462 603 1484 607
rect 29 576 37 580
rect 1024 576 1028 589
rect 29 571 1028 576
rect 1050 584 1053 585
rect 1436 584 1439 591
rect 1050 580 1441 584
rect 29 502 37 571
rect 1026 558 1041 562
rect 87 536 528 540
rect 87 514 91 536
rect 169 527 170 530
rect 385 527 578 528
rect 584 527 628 529
rect 169 526 628 527
rect 677 526 721 529
rect 764 528 808 529
rect 764 526 816 528
rect 164 525 816 526
rect 164 523 590 525
rect 164 519 188 523
rect 192 519 198 523
rect 202 519 275 523
rect 279 519 285 523
rect 289 519 368 523
rect 372 519 378 523
rect 382 522 590 523
rect 382 519 388 522
rect 584 521 590 522
rect 594 521 600 525
rect 604 522 683 525
rect 604 521 628 522
rect 677 521 683 522
rect 687 521 693 525
rect 697 522 770 525
rect 697 521 721 522
rect 764 521 770 522
rect 774 521 780 525
rect 784 522 816 525
rect 784 521 808 522
rect 168 509 169 513
rect 173 509 188 513
rect 125 502 164 505
rect 168 502 180 506
rect 29 500 89 502
rect 125 500 128 502
rect 29 497 128 500
rect 175 497 180 502
rect 184 505 188 509
rect 192 511 204 514
rect 192 508 199 511
rect 203 507 204 511
rect 255 509 256 513
rect 260 509 275 513
rect 199 506 204 507
rect 184 501 196 505
rect 192 497 196 501
rect 29 495 89 497
rect 175 493 182 497
rect 186 493 189 497
rect 168 480 172 489
rect 176 485 181 489
rect 192 482 196 493
rect 200 492 204 506
rect 256 502 267 506
rect 262 497 267 502
rect 271 505 275 509
rect 279 511 291 514
rect 279 508 286 511
rect 290 507 291 511
rect 348 509 349 513
rect 353 509 368 513
rect 286 506 291 507
rect 271 501 283 505
rect 279 497 283 501
rect 262 493 269 497
rect 273 493 276 497
rect 200 489 229 492
rect 200 488 204 489
rect 161 476 172 480
rect 179 480 196 482
rect 183 478 196 480
rect 199 487 204 488
rect 203 483 204 487
rect 199 480 204 483
rect 179 473 183 476
rect 203 476 204 480
rect 199 475 204 476
rect 168 469 169 473
rect 173 469 174 473
rect 168 463 174 469
rect 179 468 183 469
rect 188 471 189 475
rect 193 471 194 475
rect 188 463 194 471
rect 164 459 198 463
rect 202 459 208 463
rect 164 455 208 459
rect 6 448 67 450
rect 165 448 169 455
rect 225 453 229 489
rect 255 479 259 489
rect 263 485 268 489
rect 279 482 283 493
rect 287 488 291 506
rect 349 502 360 506
rect 355 497 360 502
rect 364 505 368 509
rect 372 511 384 514
rect 588 513 600 516
rect 372 508 379 511
rect 383 507 384 511
rect 397 507 466 511
rect 472 507 569 511
rect 574 507 575 511
rect 588 509 589 513
rect 593 510 600 513
rect 604 511 619 515
rect 623 511 624 515
rect 681 513 693 516
rect 588 508 593 509
rect 379 506 384 507
rect 364 501 376 505
rect 372 497 376 501
rect 355 493 362 497
rect 366 493 369 497
rect 252 476 259 479
rect 266 480 283 482
rect 270 478 283 480
rect 286 487 291 488
rect 290 483 291 487
rect 286 480 291 483
rect 266 473 270 476
rect 290 478 291 480
rect 290 476 297 478
rect 286 475 297 476
rect 348 479 352 489
rect 356 485 361 489
rect 372 482 376 493
rect 380 501 384 506
rect 380 498 474 501
rect 380 488 384 498
rect 588 501 592 508
rect 604 507 608 511
rect 681 509 682 513
rect 686 510 693 513
rect 697 511 712 515
rect 716 511 717 515
rect 768 513 780 516
rect 681 508 686 509
rect 532 497 592 501
rect 345 476 352 479
rect 359 480 376 482
rect 363 478 376 480
rect 379 487 384 488
rect 383 483 384 487
rect 397 485 454 488
rect 588 490 592 497
rect 596 503 608 507
rect 612 505 623 508
rect 596 499 600 503
rect 612 499 617 505
rect 603 495 606 499
rect 610 495 617 499
rect 681 497 685 508
rect 697 507 701 511
rect 768 509 769 513
rect 773 510 780 513
rect 784 511 799 515
rect 803 511 804 515
rect 768 508 773 509
rect 588 489 593 490
rect 460 485 570 488
rect 588 485 589 489
rect 379 480 384 483
rect 588 482 593 485
rect 255 469 256 473
rect 260 469 261 473
rect 255 463 261 469
rect 266 468 270 469
rect 275 471 276 475
rect 280 471 281 475
rect 359 473 363 476
rect 383 476 384 480
rect 379 475 384 476
rect 275 463 281 471
rect 348 469 349 473
rect 353 469 354 473
rect 348 463 354 469
rect 359 468 363 469
rect 368 471 369 475
rect 373 471 374 475
rect 534 475 556 479
rect 588 478 589 482
rect 596 484 600 495
rect 658 494 685 497
rect 611 487 616 491
rect 596 482 613 484
rect 596 480 609 482
rect 588 477 593 478
rect 620 481 624 491
rect 658 482 662 494
rect 620 478 627 481
rect 368 463 374 471
rect 435 470 439 474
rect 598 473 599 477
rect 603 473 604 477
rect 397 467 571 470
rect 598 465 604 473
rect 609 475 613 478
rect 681 490 685 494
rect 689 503 701 507
rect 705 507 719 508
rect 705 505 716 507
rect 689 499 693 503
rect 705 499 710 505
rect 696 495 699 499
rect 703 495 710 499
rect 681 489 686 490
rect 681 485 682 489
rect 681 482 686 485
rect 681 478 682 482
rect 689 484 693 495
rect 768 494 772 508
rect 784 507 788 511
rect 704 487 709 491
rect 689 482 706 484
rect 689 480 702 482
rect 681 477 686 478
rect 713 481 717 491
rect 746 490 772 494
rect 776 503 788 507
rect 792 507 806 508
rect 792 505 803 507
rect 776 499 780 503
rect 792 499 797 505
rect 1050 506 1053 580
rect 1066 573 1099 577
rect 1095 570 1099 573
rect 1152 573 1155 580
rect 1095 566 1096 570
rect 1064 558 1174 562
rect 1061 557 1174 558
rect 1450 549 1455 551
rect 1147 546 1455 549
rect 1064 525 1430 528
rect 1080 506 1083 525
rect 1125 508 1129 510
rect 807 503 1054 506
rect 1080 500 1084 502
rect 783 495 786 499
rect 790 495 797 499
rect 1014 497 1084 500
rect 713 478 720 481
rect 732 480 733 484
rect 609 470 613 471
rect 618 471 619 475
rect 623 471 624 475
rect 618 465 624 471
rect 691 473 692 477
rect 696 473 697 477
rect 691 465 697 473
rect 702 475 706 478
rect 702 470 706 471
rect 711 471 712 475
rect 716 471 717 475
rect 711 465 717 471
rect 251 459 285 463
rect 289 459 295 463
rect 251 458 295 459
rect 344 459 378 463
rect 382 459 388 463
rect 251 455 278 458
rect 344 455 388 459
rect 584 461 590 465
rect 594 461 628 465
rect 677 461 683 465
rect 687 461 721 465
rect 584 457 628 461
rect 253 448 257 455
rect 290 451 323 454
rect 344 448 348 455
rect 620 453 624 457
rect 639 456 669 459
rect 677 457 721 461
rect 732 460 736 480
rect 578 452 682 453
rect 578 450 704 452
rect 713 450 717 457
rect 746 459 750 490
rect 768 489 773 490
rect 768 485 769 489
rect 756 460 760 480
rect 768 482 773 485
rect 768 478 769 482
rect 776 484 780 495
rect 791 487 796 491
rect 776 482 793 484
rect 776 480 789 482
rect 768 477 773 478
rect 800 482 804 491
rect 800 478 808 482
rect 778 473 779 477
rect 783 473 784 477
rect 778 465 784 473
rect 789 475 793 478
rect 789 470 793 471
rect 798 471 799 475
rect 803 471 804 475
rect 798 465 804 471
rect 764 461 770 465
rect 774 461 808 465
rect 764 457 808 461
rect 802 450 806 457
rect 1014 453 1017 497
rect 1037 489 1082 492
rect 1125 491 1129 502
rect 1108 487 1111 490
rect 1125 481 1128 491
rect 1152 488 1155 512
rect 1163 506 1166 525
rect 1226 506 1229 525
rect 1236 520 1239 525
rect 1280 506 1283 525
rect 1290 520 1293 525
rect 1336 506 1339 525
rect 1346 520 1349 525
rect 1390 506 1393 525
rect 1400 520 1403 525
rect 1152 485 1176 488
rect 1180 486 1183 489
rect 1125 477 1126 481
rect 1197 480 1200 502
rect 1210 497 1213 502
rect 1243 497 1246 502
rect 1210 494 1246 497
rect 1212 486 1214 489
rect 1234 486 1235 489
rect 1243 485 1246 494
rect 1264 497 1267 502
rect 1297 497 1300 502
rect 1264 494 1300 497
rect 1320 497 1323 502
rect 1353 497 1356 502
rect 1320 494 1356 497
rect 1374 497 1377 502
rect 1407 497 1410 502
rect 1374 494 1410 497
rect 1250 485 1253 494
rect 1264 489 1271 490
rect 1264 487 1268 489
rect 1285 485 1289 488
rect 1243 482 1253 485
rect 1125 469 1128 477
rect 1197 476 1198 480
rect 1197 468 1200 476
rect 1243 469 1246 482
rect 1285 481 1288 485
rect 1297 482 1300 494
rect 1353 493 1356 494
rect 1321 486 1324 489
rect 1297 479 1316 482
rect 1297 469 1300 479
rect 1345 483 1348 485
rect 1333 475 1336 481
rect 1347 479 1348 483
rect 1345 478 1348 479
rect 1310 472 1336 475
rect 1353 469 1356 489
rect 1377 485 1378 488
rect 1396 489 1402 490
rect 1396 487 1399 489
rect 1377 476 1380 485
rect 1407 484 1410 494
rect 1379 472 1380 476
rect 1407 469 1410 480
rect 1091 459 1094 465
rect 1163 459 1166 464
rect 1209 459 1212 465
rect 1263 459 1266 465
rect 1319 459 1322 465
rect 1373 459 1376 465
rect 1055 456 1412 459
rect 1055 455 1070 456
rect 816 450 1018 453
rect 360 449 1018 450
rect 360 448 748 449
rect 6 447 283 448
rect 296 447 748 448
rect 6 446 748 447
rect 6 444 421 446
rect 6 440 92 444
rect 96 440 106 444
rect 110 440 120 444
rect 124 441 203 444
rect 124 440 187 441
rect 6 438 67 440
rect 76 439 91 440
rect 56 329 60 438
rect 90 420 94 427
rect 90 419 95 420
rect 90 415 91 419
rect 98 419 102 440
rect 105 434 118 435
rect 105 430 108 434
rect 112 430 114 434
rect 105 429 118 430
rect 105 422 111 429
rect 121 423 125 440
rect 191 440 203 441
rect 207 441 287 444
rect 207 440 271 441
rect 168 429 180 435
rect 187 434 191 437
rect 275 440 287 441
rect 291 440 324 444
rect 328 440 338 444
rect 342 440 352 444
rect 356 442 421 444
rect 425 442 435 446
rect 439 442 449 446
rect 453 443 532 446
rect 453 442 516 443
rect 356 440 391 442
rect 201 431 223 435
rect 227 431 228 435
rect 252 434 264 435
rect 201 430 205 431
rect 187 429 191 430
rect 168 426 173 429
rect 168 425 169 426
rect 98 415 101 419
rect 105 415 106 419
rect 110 415 111 419
rect 115 415 116 419
rect 121 418 125 419
rect 160 422 169 425
rect 194 426 205 430
rect 252 430 257 434
rect 261 430 264 434
rect 252 429 264 430
rect 271 434 275 437
rect 285 431 307 435
rect 311 431 312 435
rect 285 430 289 431
rect 271 429 275 430
rect 194 422 198 426
rect 212 423 213 427
rect 217 423 228 427
rect 90 414 95 415
rect 90 406 94 414
rect 110 410 116 415
rect 97 406 98 410
rect 102 406 116 410
rect 122 408 126 411
rect 160 408 163 422
rect 168 421 173 422
rect 177 420 198 422
rect 90 397 94 402
rect 90 396 95 397
rect 90 392 91 396
rect 95 392 102 395
rect 90 389 102 392
rect 106 393 110 406
rect 169 416 177 417
rect 181 418 198 420
rect 169 413 181 416
rect 122 402 126 404
rect 113 398 117 402
rect 121 398 126 402
rect 113 397 126 398
rect 169 401 173 413
rect 194 411 198 418
rect 202 416 203 420
rect 207 419 208 420
rect 207 416 219 419
rect 202 415 219 416
rect 215 412 219 415
rect 215 411 220 412
rect 183 405 189 410
rect 194 407 206 411
rect 210 407 211 411
rect 215 407 216 411
rect 183 403 185 405
rect 176 401 185 403
rect 215 406 220 407
rect 224 407 228 423
rect 252 426 257 429
rect 252 422 253 426
rect 278 426 289 430
rect 278 422 282 426
rect 296 423 297 427
rect 301 423 312 427
rect 252 421 257 422
rect 261 420 282 422
rect 253 416 261 417
rect 265 418 282 420
rect 253 413 265 416
rect 215 402 219 406
rect 176 397 189 401
rect 195 398 219 402
rect 224 403 226 407
rect 169 396 173 397
rect 195 396 199 398
rect 106 389 120 393
rect 124 389 125 393
rect 182 389 183 393
rect 187 389 188 393
rect 224 394 228 403
rect 253 401 257 413
rect 278 411 282 418
rect 286 416 287 420
rect 291 419 292 420
rect 291 416 303 419
rect 286 415 303 416
rect 299 412 303 415
rect 308 414 312 423
rect 322 420 326 427
rect 322 419 327 420
rect 322 415 323 419
rect 330 419 334 440
rect 337 434 346 435
rect 337 430 340 434
rect 344 431 346 434
rect 344 430 350 431
rect 337 429 350 430
rect 337 422 343 429
rect 353 423 357 440
rect 364 423 382 426
rect 330 415 333 419
rect 337 415 338 419
rect 342 415 343 419
rect 347 415 348 419
rect 353 418 357 419
rect 299 411 304 412
rect 267 405 273 410
rect 278 407 290 411
rect 294 407 295 411
rect 299 407 300 411
rect 267 403 269 405
rect 260 401 269 403
rect 299 406 304 407
rect 308 411 315 414
rect 322 414 327 415
rect 299 402 303 406
rect 260 397 273 401
rect 279 398 303 402
rect 253 396 257 397
rect 279 396 283 398
rect 195 391 199 392
rect 204 390 205 394
rect 209 390 228 394
rect 182 384 188 389
rect 266 389 267 393
rect 271 389 272 393
rect 308 394 312 411
rect 322 406 326 414
rect 342 410 348 415
rect 329 406 330 410
rect 334 406 348 410
rect 354 409 358 411
rect 279 391 283 392
rect 288 390 289 394
rect 293 390 312 394
rect 316 403 326 406
rect 316 391 319 403
rect 266 384 272 389
rect 322 397 326 403
rect 322 396 327 397
rect 322 392 323 396
rect 327 392 334 395
rect 322 389 334 392
rect 338 393 342 406
rect 354 402 358 405
rect 345 398 349 402
rect 353 398 358 402
rect 345 397 358 398
rect 338 389 352 393
rect 356 389 357 393
rect 89 380 92 384
rect 96 380 102 384
rect 106 380 170 384
rect 174 380 223 384
rect 227 380 254 384
rect 258 380 307 384
rect 311 380 324 384
rect 328 380 334 384
rect 338 383 362 384
rect 338 380 356 383
rect 75 377 356 380
rect 75 376 362 377
rect 179 374 223 376
rect 179 370 185 374
rect 189 370 213 374
rect 217 370 223 374
rect 183 362 189 370
rect 183 358 184 362
rect 188 358 189 362
rect 194 362 198 363
rect 203 362 209 370
rect 203 358 204 362
rect 208 358 209 362
rect 214 362 219 365
rect 377 366 381 423
rect 350 363 382 366
rect 218 358 219 362
rect 194 355 198 358
rect 214 357 219 358
rect 194 351 211 355
rect 183 339 187 349
rect 191 344 196 348
rect 207 347 211 351
rect 191 336 197 340
rect 201 336 204 340
rect 55 309 60 329
rect 191 330 195 336
rect 207 332 211 343
rect 178 327 195 330
rect 199 328 211 332
rect 215 353 376 357
rect 199 324 203 328
rect 215 327 219 353
rect 385 331 389 440
rect 419 422 423 429
rect 419 421 424 422
rect 419 417 420 421
rect 427 421 431 442
rect 434 436 447 437
rect 434 432 437 436
rect 441 432 443 436
rect 434 431 447 432
rect 434 424 440 431
rect 450 425 454 442
rect 520 442 532 443
rect 536 443 616 446
rect 536 442 600 443
rect 497 431 509 437
rect 516 436 520 439
rect 604 442 616 443
rect 620 442 653 446
rect 657 442 667 446
rect 671 442 681 446
rect 685 445 748 446
rect 752 445 762 449
rect 766 445 776 449
rect 780 446 859 449
rect 780 445 843 446
rect 685 442 721 445
rect 530 433 552 437
rect 556 433 557 437
rect 572 436 593 437
rect 530 432 534 433
rect 516 431 520 432
rect 497 428 502 431
rect 497 427 498 428
rect 427 417 430 421
rect 434 417 435 421
rect 439 417 440 421
rect 444 417 445 421
rect 450 420 454 421
rect 489 424 498 427
rect 523 428 534 432
rect 572 432 586 436
rect 590 432 593 436
rect 572 431 593 432
rect 600 436 604 439
rect 614 433 636 437
rect 640 433 641 437
rect 614 432 618 433
rect 600 431 604 432
rect 523 424 527 428
rect 541 425 542 429
rect 546 425 557 429
rect 419 416 424 417
rect 419 408 423 416
rect 439 412 445 417
rect 426 408 427 412
rect 431 408 445 412
rect 451 410 455 413
rect 489 410 492 424
rect 497 423 502 424
rect 506 422 527 424
rect 419 399 423 404
rect 419 398 424 399
rect 419 394 420 398
rect 424 394 431 397
rect 419 391 431 394
rect 435 395 439 408
rect 498 418 506 419
rect 510 420 527 422
rect 498 415 510 418
rect 451 404 455 406
rect 442 400 446 404
rect 450 400 455 404
rect 442 399 455 400
rect 498 403 502 415
rect 523 413 527 420
rect 531 418 532 422
rect 536 421 537 422
rect 536 418 548 421
rect 531 417 548 418
rect 544 414 548 417
rect 544 413 549 414
rect 512 407 518 412
rect 523 409 535 413
rect 539 409 540 413
rect 544 409 545 413
rect 512 405 514 407
rect 505 403 514 405
rect 544 408 549 409
rect 553 409 557 425
rect 581 428 586 431
rect 581 424 582 428
rect 607 428 618 432
rect 607 424 611 428
rect 625 425 626 429
rect 630 425 643 429
rect 581 423 586 424
rect 590 422 611 424
rect 582 418 590 419
rect 594 420 611 422
rect 582 415 594 418
rect 544 404 548 408
rect 505 399 518 403
rect 524 400 548 404
rect 553 405 555 409
rect 498 398 502 399
rect 524 398 528 400
rect 435 391 449 395
rect 453 391 454 395
rect 511 391 512 395
rect 516 391 517 395
rect 553 396 557 405
rect 582 403 586 415
rect 607 413 611 420
rect 615 418 616 422
rect 620 421 621 422
rect 620 418 632 421
rect 615 417 632 418
rect 628 414 632 417
rect 628 413 633 414
rect 596 407 602 412
rect 607 409 619 413
rect 623 409 624 413
rect 628 409 629 413
rect 596 405 598 407
rect 589 403 598 405
rect 628 408 633 409
rect 628 404 632 408
rect 589 399 602 403
rect 608 400 632 404
rect 582 398 586 399
rect 608 398 612 400
rect 524 393 528 394
rect 533 392 534 396
rect 538 392 557 396
rect 511 386 517 391
rect 595 391 596 395
rect 600 391 601 395
rect 637 396 641 425
rect 651 422 655 429
rect 651 421 656 422
rect 651 417 652 421
rect 659 421 663 442
rect 666 436 679 437
rect 666 432 669 436
rect 673 432 675 436
rect 666 431 679 432
rect 666 424 672 431
rect 682 425 686 442
rect 659 417 662 421
rect 666 417 667 421
rect 671 417 672 421
rect 676 417 677 421
rect 682 420 686 421
rect 651 416 656 417
rect 651 408 655 416
rect 671 412 677 417
rect 658 408 659 412
rect 663 408 677 412
rect 683 411 687 413
rect 608 393 612 394
rect 617 392 618 396
rect 622 392 641 396
rect 645 405 655 408
rect 645 393 648 405
rect 595 386 601 391
rect 651 399 655 405
rect 651 398 656 399
rect 651 394 652 398
rect 656 394 663 397
rect 651 391 663 394
rect 667 395 671 408
rect 683 404 687 407
rect 674 400 678 404
rect 682 400 687 404
rect 674 399 687 400
rect 667 391 681 395
rect 685 391 686 395
rect 418 382 421 386
rect 425 382 431 386
rect 435 382 499 386
rect 503 382 552 386
rect 556 382 583 386
rect 587 382 636 386
rect 640 382 653 386
rect 657 382 663 386
rect 667 385 691 386
rect 667 382 683 385
rect 418 381 683 382
rect 403 379 683 381
rect 689 379 691 385
rect 403 378 691 379
rect 403 377 419 378
rect 508 376 552 378
rect 508 372 514 376
rect 518 372 542 376
rect 546 372 552 376
rect 405 353 473 357
rect 214 326 219 327
rect 183 320 184 324
rect 188 320 203 324
rect 206 322 214 324
rect 218 322 219 326
rect 349 325 376 329
rect 206 320 219 322
rect 201 314 202 317
rect 179 313 202 314
rect 206 314 207 317
rect 206 313 213 314
rect 179 310 213 313
rect 217 310 223 314
rect 179 309 223 310
rect 384 311 389 331
rect 487 330 490 365
rect 512 364 518 372
rect 512 360 513 364
rect 517 360 518 364
rect 523 364 527 365
rect 532 364 538 372
rect 532 360 533 364
rect 537 360 538 364
rect 543 364 548 367
rect 588 365 672 368
rect 547 360 548 364
rect 523 357 527 360
rect 543 359 548 360
rect 523 353 540 357
rect 512 341 516 351
rect 520 346 525 350
rect 536 349 540 353
rect 520 338 526 342
rect 530 338 533 342
rect 520 332 524 338
rect 536 334 540 345
rect 507 329 524 332
rect 528 330 540 334
rect 544 353 548 359
rect 544 350 695 353
rect 699 350 700 353
rect 528 326 532 330
rect 544 329 548 350
rect 712 334 716 442
rect 746 425 750 432
rect 746 424 751 425
rect 746 420 747 424
rect 754 424 758 445
rect 761 439 774 440
rect 761 435 764 439
rect 768 435 770 439
rect 761 434 774 435
rect 761 427 767 434
rect 777 428 781 445
rect 847 445 859 446
rect 863 446 943 449
rect 863 445 927 446
rect 824 434 836 440
rect 843 439 847 442
rect 931 445 943 446
rect 947 445 980 449
rect 984 445 994 449
rect 998 445 1008 449
rect 1012 445 1018 449
rect 857 436 879 440
rect 883 436 884 440
rect 897 439 920 440
rect 857 435 861 436
rect 897 435 913 439
rect 917 435 920 439
rect 843 434 847 435
rect 824 431 829 434
rect 824 430 825 431
rect 754 420 757 424
rect 761 420 762 424
rect 766 420 767 424
rect 771 420 772 424
rect 777 423 781 424
rect 746 419 751 420
rect 746 411 750 419
rect 766 415 772 420
rect 753 411 754 415
rect 758 411 772 415
rect 778 413 782 416
rect 746 402 750 407
rect 746 401 751 402
rect 746 397 747 401
rect 751 397 758 400
rect 746 394 758 397
rect 762 398 766 411
rect 778 407 782 409
rect 769 403 773 407
rect 777 403 782 407
rect 769 402 782 403
rect 791 398 794 417
rect 762 394 776 398
rect 780 394 781 398
rect 792 394 794 398
rect 805 396 809 425
rect 816 427 825 430
rect 850 431 861 435
rect 850 427 854 431
rect 868 428 869 432
rect 873 428 884 432
rect 816 413 819 427
rect 824 426 829 427
rect 833 425 854 427
rect 825 421 833 422
rect 837 423 854 425
rect 825 418 837 421
rect 825 406 829 418
rect 850 416 854 423
rect 858 421 859 425
rect 863 424 864 425
rect 863 421 875 424
rect 858 420 875 421
rect 871 417 875 420
rect 871 416 876 417
rect 839 410 845 415
rect 850 412 862 416
rect 866 412 867 416
rect 871 412 872 416
rect 839 408 841 410
rect 832 406 841 408
rect 871 411 876 412
rect 880 412 884 428
rect 871 407 875 411
rect 832 402 845 406
rect 851 403 875 407
rect 880 408 882 412
rect 825 401 829 402
rect 851 401 855 403
rect 805 392 806 396
rect 838 394 839 398
rect 843 394 844 398
rect 880 399 884 408
rect 851 396 855 397
rect 860 395 861 399
rect 865 395 884 399
rect 891 396 894 427
rect 838 389 844 394
rect 898 389 902 435
rect 908 434 920 435
rect 927 439 931 442
rect 941 436 963 440
rect 967 436 968 440
rect 941 435 945 436
rect 927 434 931 435
rect 908 431 913 434
rect 908 427 909 431
rect 934 431 945 435
rect 934 427 938 431
rect 952 428 953 432
rect 957 428 968 432
rect 908 426 913 427
rect 917 425 938 427
rect 909 421 917 422
rect 921 423 938 425
rect 909 418 921 421
rect 909 406 913 418
rect 934 416 938 423
rect 942 421 943 425
rect 947 424 948 425
rect 947 421 959 424
rect 942 420 959 421
rect 955 417 959 420
rect 955 416 960 417
rect 923 410 929 415
rect 934 412 946 416
rect 950 412 951 416
rect 955 412 956 416
rect 923 408 925 410
rect 916 406 925 408
rect 955 411 960 412
rect 955 407 959 411
rect 916 402 929 406
rect 935 403 959 407
rect 909 401 913 402
rect 935 401 939 403
rect 922 394 923 398
rect 927 394 928 398
rect 964 399 968 428
rect 978 425 982 432
rect 978 424 983 425
rect 978 420 979 424
rect 986 424 990 445
rect 993 439 1006 440
rect 993 435 996 439
rect 1000 435 1002 439
rect 993 434 1006 435
rect 993 427 999 434
rect 1009 428 1013 445
rect 986 420 989 424
rect 993 420 994 424
rect 998 420 999 424
rect 1003 420 1004 424
rect 1009 423 1013 424
rect 978 419 983 420
rect 978 411 982 419
rect 998 415 1004 420
rect 985 411 986 415
rect 990 411 1004 415
rect 1010 414 1014 416
rect 935 396 939 397
rect 944 395 945 399
rect 949 395 968 399
rect 972 408 982 411
rect 972 396 975 408
rect 922 389 928 394
rect 978 402 982 408
rect 978 401 983 402
rect 978 397 979 401
rect 983 397 990 400
rect 978 394 990 397
rect 994 398 998 411
rect 1010 407 1014 410
rect 1001 403 1005 407
rect 1009 403 1014 407
rect 1001 402 1014 403
rect 994 394 1008 398
rect 1012 394 1013 398
rect 745 388 748 389
rect 743 385 748 388
rect 752 385 758 389
rect 762 385 826 389
rect 830 385 879 389
rect 883 385 910 389
rect 914 385 963 389
rect 967 385 980 389
rect 984 385 990 389
rect 994 385 1018 389
rect 743 383 1018 385
rect 730 381 1018 383
rect 730 380 747 381
rect 730 379 746 380
rect 835 379 879 381
rect 835 375 841 379
rect 845 375 869 379
rect 873 375 879 379
rect 839 367 845 375
rect 543 328 548 329
rect 512 322 513 326
rect 517 322 532 326
rect 535 324 543 326
rect 547 324 548 328
rect 535 322 548 324
rect 673 319 676 333
rect 530 316 531 319
rect 508 315 531 316
rect 535 316 536 319
rect 673 316 702 319
rect 535 315 542 316
rect 508 312 542 315
rect 546 312 552 316
rect 508 311 552 312
rect 55 306 223 309
rect 55 305 183 306
rect 361 305 376 309
rect 180 302 183 305
rect 384 308 552 311
rect 384 307 510 308
rect 507 304 510 307
rect 55 298 361 302
rect 55 294 91 298
rect 95 294 105 298
rect 109 294 119 298
rect 123 295 202 298
rect 123 294 186 295
rect 55 183 59 294
rect 89 274 93 281
rect 89 273 94 274
rect 89 269 90 273
rect 97 273 101 294
rect 104 288 117 289
rect 104 284 107 288
rect 111 284 113 288
rect 104 283 117 284
rect 104 276 110 283
rect 120 277 124 294
rect 190 294 202 295
rect 206 295 286 298
rect 206 294 270 295
rect 167 283 179 289
rect 186 288 190 291
rect 274 294 286 295
rect 290 294 323 298
rect 327 294 337 298
rect 341 294 351 298
rect 355 294 361 298
rect 384 300 690 304
rect 384 296 420 300
rect 424 296 434 300
rect 438 296 448 300
rect 452 297 531 300
rect 452 296 515 297
rect 200 285 222 289
rect 226 285 227 289
rect 251 288 263 289
rect 239 285 256 288
rect 200 284 204 285
rect 186 283 190 284
rect 167 280 172 283
rect 167 279 168 280
rect 97 269 100 273
rect 104 269 105 273
rect 109 269 110 273
rect 114 269 115 273
rect 120 272 124 273
rect 159 276 168 279
rect 193 280 204 284
rect 193 276 197 280
rect 211 277 212 281
rect 216 277 227 281
rect 89 268 94 269
rect 89 260 93 268
rect 109 264 115 269
rect 96 260 97 264
rect 101 260 115 264
rect 121 262 125 265
rect 159 262 162 276
rect 167 275 172 276
rect 176 274 197 276
rect 89 251 93 256
rect 89 250 94 251
rect 89 246 90 250
rect 94 246 101 249
rect 89 243 101 246
rect 105 247 109 260
rect 168 270 176 271
rect 180 272 197 274
rect 168 267 180 270
rect 121 256 125 258
rect 112 252 116 256
rect 120 252 125 256
rect 112 251 125 252
rect 168 255 172 267
rect 193 265 197 272
rect 201 270 202 274
rect 206 273 207 274
rect 206 270 218 273
rect 201 269 218 270
rect 214 266 218 269
rect 214 265 219 266
rect 182 259 188 264
rect 193 261 205 265
rect 209 261 210 265
rect 214 261 215 265
rect 182 257 184 259
rect 175 255 184 257
rect 214 260 219 261
rect 223 261 227 277
rect 214 256 218 260
rect 175 251 188 255
rect 194 252 218 256
rect 223 257 225 261
rect 168 250 172 251
rect 194 250 198 252
rect 105 243 119 247
rect 123 243 124 247
rect 181 243 182 247
rect 186 243 187 247
rect 223 248 227 257
rect 194 245 198 246
rect 203 244 204 248
rect 208 244 227 248
rect 239 245 242 285
rect 251 284 256 285
rect 260 284 263 288
rect 251 283 263 284
rect 270 288 274 291
rect 284 285 306 289
rect 310 285 311 289
rect 284 284 288 285
rect 270 283 274 284
rect 251 280 256 283
rect 251 276 252 280
rect 277 280 288 284
rect 277 276 281 280
rect 295 277 296 281
rect 300 277 311 281
rect 251 275 256 276
rect 260 274 281 276
rect 307 275 311 277
rect 252 270 260 271
rect 264 272 281 274
rect 252 267 264 270
rect 252 255 256 267
rect 277 265 281 272
rect 285 270 286 274
rect 290 273 291 274
rect 290 270 302 273
rect 285 269 302 270
rect 298 266 302 269
rect 307 272 314 275
rect 321 274 325 281
rect 321 273 326 274
rect 298 265 303 266
rect 266 259 272 264
rect 277 261 289 265
rect 293 261 294 265
rect 298 261 299 265
rect 266 257 268 259
rect 259 255 268 257
rect 298 260 303 261
rect 298 256 302 260
rect 259 251 272 255
rect 278 252 302 256
rect 252 250 256 251
rect 278 250 282 252
rect 181 238 187 243
rect 265 243 266 247
rect 270 243 271 247
rect 307 248 311 272
rect 321 269 322 273
rect 329 273 333 294
rect 336 288 349 289
rect 336 284 339 288
rect 343 284 345 288
rect 336 283 349 284
rect 336 276 342 283
rect 352 277 356 294
rect 365 276 376 279
rect 329 269 332 273
rect 336 269 337 273
rect 341 269 342 273
rect 346 269 347 273
rect 352 272 356 273
rect 321 268 326 269
rect 321 260 325 268
rect 341 264 347 269
rect 328 260 329 264
rect 333 260 347 264
rect 353 263 357 265
rect 278 245 282 246
rect 287 244 288 248
rect 292 244 311 248
rect 315 257 325 260
rect 315 245 318 257
rect 265 238 271 243
rect 321 251 325 257
rect 321 250 326 251
rect 321 246 322 250
rect 326 246 333 249
rect 321 243 333 246
rect 337 247 341 260
rect 353 256 357 259
rect 344 252 348 256
rect 352 252 357 256
rect 344 251 357 252
rect 337 243 351 247
rect 355 243 356 247
rect 88 234 91 238
rect 95 234 101 238
rect 105 234 169 238
rect 173 234 222 238
rect 226 234 253 238
rect 257 234 306 238
rect 310 234 323 238
rect 327 234 333 238
rect 337 234 356 238
rect 88 231 356 234
rect 88 230 361 231
rect 178 228 222 230
rect 178 224 184 228
rect 188 224 212 228
rect 216 224 222 228
rect 182 216 188 224
rect 182 212 183 216
rect 187 212 188 216
rect 193 216 197 217
rect 202 216 208 224
rect 309 221 350 224
rect 202 212 203 216
rect 207 212 208 216
rect 213 216 218 219
rect 217 212 218 216
rect 193 209 197 212
rect 213 211 218 212
rect 193 205 210 209
rect 182 193 186 203
rect 190 198 195 202
rect 206 201 210 205
rect 190 190 196 194
rect 200 190 203 194
rect 54 163 59 183
rect 190 184 194 190
rect 206 186 210 197
rect 177 181 194 184
rect 198 182 210 186
rect 214 199 218 211
rect 306 203 329 206
rect 334 203 335 206
rect 214 196 293 199
rect 198 178 202 182
rect 214 181 218 196
rect 213 180 218 181
rect 182 174 183 178
rect 187 174 202 178
rect 205 176 213 178
rect 217 176 218 180
rect 290 181 293 196
rect 290 178 336 181
rect 205 174 218 176
rect 200 168 201 171
rect 178 167 201 168
rect 205 168 206 171
rect 205 167 212 168
rect 178 164 212 167
rect 216 164 222 168
rect 178 163 222 164
rect 54 160 222 163
rect 54 159 178 160
rect 347 120 350 221
rect 359 202 375 206
rect 384 185 388 296
rect 418 276 422 283
rect 418 275 423 276
rect 418 271 419 275
rect 426 275 430 296
rect 433 290 446 291
rect 433 286 436 290
rect 440 286 442 290
rect 433 285 446 286
rect 433 278 439 285
rect 449 279 453 296
rect 519 296 531 297
rect 535 297 615 300
rect 535 296 599 297
rect 496 285 508 291
rect 515 290 519 293
rect 603 296 615 297
rect 619 296 652 300
rect 656 296 666 300
rect 670 296 680 300
rect 684 296 690 300
rect 529 287 551 291
rect 555 287 556 291
rect 580 290 592 291
rect 529 286 533 287
rect 515 285 519 286
rect 496 282 501 285
rect 496 281 497 282
rect 426 271 429 275
rect 433 271 434 275
rect 438 271 439 275
rect 443 271 444 275
rect 449 274 453 275
rect 488 278 497 281
rect 522 282 533 286
rect 580 286 585 290
rect 589 286 592 290
rect 580 285 592 286
rect 599 290 603 293
rect 613 287 635 291
rect 639 287 640 291
rect 613 286 617 287
rect 599 285 603 286
rect 522 278 526 282
rect 540 279 541 283
rect 545 279 556 283
rect 418 270 423 271
rect 418 262 422 270
rect 438 266 444 271
rect 425 262 426 266
rect 430 262 444 266
rect 450 264 454 267
rect 418 253 422 258
rect 418 252 423 253
rect 418 248 419 252
rect 423 248 430 251
rect 418 245 430 248
rect 434 249 438 262
rect 450 258 454 260
rect 441 254 445 258
rect 449 254 454 258
rect 441 253 454 254
rect 434 245 448 249
rect 452 245 453 249
rect 478 247 481 267
rect 488 264 491 278
rect 496 277 501 278
rect 505 276 526 278
rect 497 272 505 273
rect 509 274 526 276
rect 497 269 509 272
rect 497 257 501 269
rect 522 267 526 274
rect 530 272 531 276
rect 535 275 536 276
rect 535 272 547 275
rect 530 271 547 272
rect 543 268 547 271
rect 543 267 548 268
rect 511 261 517 266
rect 522 263 534 267
rect 538 263 539 267
rect 543 263 544 267
rect 511 259 513 261
rect 504 257 513 259
rect 543 262 548 263
rect 552 263 556 279
rect 580 282 585 285
rect 580 278 581 282
rect 606 282 617 286
rect 606 278 610 282
rect 624 279 625 283
rect 629 279 640 283
rect 580 277 585 278
rect 589 276 610 278
rect 581 272 589 273
rect 593 274 610 276
rect 581 269 593 272
rect 543 258 547 262
rect 504 253 517 257
rect 523 254 547 258
rect 552 259 554 263
rect 497 252 501 253
rect 523 252 527 254
rect 510 245 511 249
rect 515 245 516 249
rect 552 250 556 259
rect 581 257 585 269
rect 606 267 610 274
rect 614 272 615 276
rect 619 275 620 276
rect 619 272 631 275
rect 614 271 631 272
rect 627 268 631 271
rect 636 273 640 279
rect 650 276 654 283
rect 650 275 655 276
rect 636 270 643 273
rect 650 271 651 275
rect 658 275 662 296
rect 665 290 678 291
rect 665 286 668 290
rect 672 286 674 290
rect 665 285 678 286
rect 665 278 671 285
rect 681 279 685 296
rect 658 271 661 275
rect 665 271 666 275
rect 670 271 671 275
rect 675 271 676 275
rect 681 274 685 275
rect 650 270 655 271
rect 627 267 632 268
rect 595 261 601 266
rect 606 263 618 267
rect 622 263 623 267
rect 627 263 628 267
rect 595 259 597 261
rect 588 257 597 259
rect 627 262 632 263
rect 627 258 631 262
rect 588 253 601 257
rect 607 254 631 258
rect 581 252 585 253
rect 607 252 611 254
rect 523 247 527 248
rect 532 246 533 250
rect 537 246 556 250
rect 510 240 516 245
rect 594 245 595 249
rect 599 245 600 249
rect 636 250 640 270
rect 650 262 654 270
rect 670 266 676 271
rect 657 262 658 266
rect 662 262 676 266
rect 682 265 686 267
rect 607 247 611 248
rect 616 246 617 250
rect 621 246 640 250
rect 644 259 654 262
rect 644 247 647 259
rect 594 240 600 245
rect 650 253 654 259
rect 650 252 655 253
rect 650 248 651 252
rect 655 248 662 251
rect 650 245 662 248
rect 666 249 670 262
rect 682 258 686 261
rect 673 254 677 258
rect 681 254 686 258
rect 673 253 686 254
rect 666 245 680 249
rect 684 245 685 249
rect 417 236 420 240
rect 424 236 430 240
rect 434 236 498 240
rect 502 236 551 240
rect 555 236 582 240
rect 586 236 635 240
rect 639 236 652 240
rect 656 236 662 240
rect 666 236 690 240
rect 398 233 683 236
rect 417 232 683 233
rect 687 232 690 236
rect 507 230 551 232
rect 427 228 489 229
rect 431 226 489 228
rect 431 225 467 226
rect 507 226 513 230
rect 517 226 541 230
rect 545 226 551 230
rect 478 221 481 223
rect 511 218 517 226
rect 406 210 454 213
rect 478 203 481 217
rect 511 214 512 218
rect 516 214 517 218
rect 522 218 526 219
rect 531 218 537 226
rect 677 228 681 229
rect 635 225 681 228
rect 531 214 532 218
rect 536 214 537 218
rect 542 218 547 221
rect 546 214 547 218
rect 522 211 526 214
rect 542 213 547 214
rect 522 207 539 211
rect 360 178 375 181
rect 383 165 388 185
rect 428 173 432 201
rect 450 199 478 202
rect 450 173 454 199
rect 511 195 515 205
rect 519 200 524 204
rect 535 203 539 207
rect 519 192 525 196
rect 529 192 532 196
rect 519 186 523 192
rect 535 188 539 199
rect 506 183 523 186
rect 527 184 539 188
rect 527 180 531 184
rect 543 183 547 213
rect 574 209 656 214
rect 677 194 681 225
rect 680 191 681 194
rect 542 182 547 183
rect 511 176 512 180
rect 516 176 531 180
rect 534 178 542 180
rect 546 180 547 182
rect 546 178 551 180
rect 534 176 551 178
rect 529 170 530 173
rect 507 169 530 170
rect 534 170 535 173
rect 534 169 541 170
rect 507 166 541 169
rect 545 166 551 170
rect 507 165 551 166
rect 383 162 551 165
rect 383 161 507 162
rect 496 154 500 161
rect 379 152 423 154
rect 472 152 516 154
rect 559 152 603 154
rect 379 150 603 152
rect 379 146 385 150
rect 389 149 478 150
rect 389 146 423 149
rect 472 146 478 149
rect 482 149 565 150
rect 482 146 516 149
rect 559 146 565 149
rect 569 146 603 150
rect 699 146 702 316
rect 711 314 716 334
rect 720 362 723 363
rect 720 359 755 362
rect 839 363 840 367
rect 844 363 845 367
rect 850 367 854 368
rect 859 367 865 375
rect 859 363 860 367
rect 864 363 865 367
rect 870 367 875 370
rect 874 363 875 367
rect 720 322 723 359
rect 731 350 798 353
rect 802 350 803 353
rect 808 322 812 362
rect 850 360 854 363
rect 870 362 875 363
rect 850 356 867 360
rect 820 328 823 355
rect 839 344 843 354
rect 847 349 852 353
rect 863 352 867 356
rect 847 341 853 345
rect 857 341 860 345
rect 847 335 851 341
rect 863 337 867 348
rect 834 332 851 335
rect 855 333 867 337
rect 871 358 875 362
rect 871 355 883 358
rect 855 329 859 333
rect 871 332 875 355
rect 1011 353 1014 381
rect 1055 353 1058 455
rect 1235 453 1240 456
rect 1341 453 1345 456
rect 1167 450 1416 453
rect 1167 445 1170 450
rect 1213 444 1216 450
rect 1267 444 1270 450
rect 1323 444 1326 450
rect 1377 444 1380 450
rect 1064 398 1068 437
rect 1201 433 1204 441
rect 1201 429 1202 433
rect 1184 420 1187 423
rect 1201 407 1204 429
rect 1247 427 1250 440
rect 1247 424 1257 427
rect 1289 424 1292 428
rect 1301 430 1304 440
rect 1301 427 1320 430
rect 1349 430 1352 431
rect 1216 420 1218 423
rect 1238 420 1239 423
rect 1247 415 1250 424
rect 1214 412 1250 415
rect 1214 407 1217 412
rect 1247 407 1250 412
rect 1254 415 1257 424
rect 1268 420 1272 422
rect 1289 421 1293 424
rect 1268 419 1275 420
rect 1301 415 1304 427
rect 1351 426 1352 430
rect 1349 424 1352 426
rect 1325 420 1328 423
rect 1357 420 1360 440
rect 1383 433 1384 437
rect 1381 424 1384 433
rect 1411 429 1414 440
rect 1381 421 1382 424
rect 1400 420 1403 422
rect 1400 419 1406 420
rect 1357 415 1360 416
rect 1411 415 1414 425
rect 1268 412 1304 415
rect 1268 407 1271 412
rect 1301 407 1304 412
rect 1324 412 1360 415
rect 1324 407 1327 412
rect 1357 407 1360 412
rect 1378 412 1414 415
rect 1378 407 1381 412
rect 1411 407 1414 412
rect 1167 384 1170 403
rect 1230 384 1233 403
rect 1240 384 1243 389
rect 1284 384 1287 403
rect 1294 384 1297 389
rect 1340 384 1343 403
rect 1350 384 1353 389
rect 1394 384 1397 403
rect 1404 384 1407 389
rect 1425 384 1430 525
rect 1450 443 1455 546
rect 1165 383 1430 384
rect 1062 381 1430 383
rect 1062 380 1428 381
rect 1078 361 1081 380
rect 1123 363 1127 365
rect 1161 361 1164 380
rect 1175 372 1204 375
rect 1011 350 1058 353
rect 891 334 894 349
rect 870 331 875 332
rect 839 325 840 329
rect 844 325 859 329
rect 862 327 870 329
rect 874 327 875 331
rect 862 325 875 327
rect 720 321 729 322
rect 720 317 739 321
rect 743 317 748 321
rect 857 319 858 322
rect 808 317 812 318
rect 835 318 858 319
rect 862 319 863 322
rect 890 321 895 334
rect 862 318 869 319
rect 835 315 869 318
rect 873 315 879 319
rect 835 314 879 315
rect 1040 317 1044 318
rect 711 311 879 314
rect 1007 314 1045 317
rect 1055 314 1058 350
rect 1123 346 1127 357
rect 1106 342 1109 345
rect 1123 336 1126 346
rect 1178 341 1181 344
rect 1123 332 1124 336
rect 1195 335 1198 357
rect 1201 345 1204 372
rect 1224 361 1227 380
rect 1234 375 1237 380
rect 1278 361 1281 380
rect 1288 375 1291 380
rect 1334 361 1337 380
rect 1344 375 1347 380
rect 1388 361 1391 380
rect 1398 375 1401 380
rect 1208 352 1211 357
rect 1241 352 1244 357
rect 1208 349 1244 352
rect 1201 342 1206 345
rect 1210 341 1212 344
rect 1232 341 1233 344
rect 1241 340 1244 349
rect 1262 352 1265 357
rect 1295 352 1298 357
rect 1262 349 1298 352
rect 1318 352 1321 357
rect 1351 352 1354 357
rect 1318 349 1354 352
rect 1372 352 1375 357
rect 1405 352 1408 357
rect 1372 349 1408 352
rect 1248 340 1251 349
rect 1262 344 1269 345
rect 1262 342 1266 344
rect 1283 340 1287 343
rect 1241 337 1251 340
rect 1123 324 1126 332
rect 1195 331 1196 335
rect 1195 323 1198 331
rect 1241 324 1244 337
rect 1283 336 1286 340
rect 1295 337 1298 349
rect 1351 348 1354 349
rect 1319 341 1322 344
rect 1295 334 1314 337
rect 1295 324 1298 334
rect 1343 338 1346 340
rect 1331 330 1334 336
rect 1345 334 1346 338
rect 1343 333 1346 334
rect 1308 327 1334 330
rect 1351 324 1354 344
rect 1375 340 1376 343
rect 1394 344 1400 345
rect 1394 342 1397 344
rect 1375 331 1378 340
rect 1405 339 1408 349
rect 1377 327 1378 331
rect 1405 324 1408 335
rect 1089 314 1092 320
rect 1161 314 1164 319
rect 1207 314 1210 320
rect 1261 314 1264 320
rect 1317 314 1320 320
rect 1371 314 1374 320
rect 711 310 835 311
rect 840 307 843 311
rect 711 303 1017 307
rect 711 299 747 303
rect 751 299 761 303
rect 765 299 775 303
rect 779 300 858 303
rect 779 299 842 300
rect 711 188 715 299
rect 745 279 749 286
rect 745 278 750 279
rect 745 274 746 278
rect 753 278 757 299
rect 760 293 773 294
rect 760 289 763 293
rect 767 289 769 293
rect 760 288 773 289
rect 760 281 766 288
rect 776 282 780 299
rect 846 299 858 300
rect 862 300 942 303
rect 862 299 926 300
rect 823 288 835 294
rect 842 293 846 296
rect 930 299 942 300
rect 946 299 979 303
rect 983 299 993 303
rect 997 299 1007 303
rect 1011 299 1017 303
rect 856 290 878 294
rect 882 290 883 294
rect 907 293 919 294
rect 856 289 860 290
rect 842 288 846 289
rect 823 285 828 288
rect 753 274 756 278
rect 760 274 761 278
rect 765 274 766 278
rect 770 274 771 278
rect 776 277 780 278
rect 823 284 824 285
rect 745 273 750 274
rect 745 265 749 273
rect 765 269 771 274
rect 752 265 753 269
rect 757 265 771 269
rect 777 267 781 270
rect 745 256 749 261
rect 745 255 750 256
rect 745 251 746 255
rect 750 251 757 254
rect 745 248 757 251
rect 761 252 765 265
rect 777 261 781 263
rect 768 257 772 261
rect 776 257 781 261
rect 768 256 781 257
rect 794 255 798 280
rect 815 281 824 284
rect 849 285 860 289
rect 907 289 912 293
rect 916 289 919 293
rect 907 288 919 289
rect 926 293 930 296
rect 940 290 962 294
rect 966 290 967 294
rect 940 289 944 290
rect 926 288 930 289
rect 849 281 853 285
rect 867 282 868 286
rect 872 282 883 286
rect 815 267 818 281
rect 823 280 828 281
rect 832 279 853 281
rect 824 275 832 276
rect 836 277 853 279
rect 824 272 836 275
rect 824 260 828 272
rect 849 270 853 277
rect 857 275 858 279
rect 862 278 863 279
rect 862 275 874 278
rect 857 274 874 275
rect 870 271 874 274
rect 870 270 875 271
rect 838 264 844 269
rect 849 266 861 270
rect 865 266 866 270
rect 870 266 871 270
rect 838 262 840 264
rect 824 255 828 256
rect 831 260 840 262
rect 870 265 875 266
rect 879 266 883 282
rect 907 285 912 288
rect 907 281 908 285
rect 933 285 944 289
rect 933 281 937 285
rect 951 282 952 286
rect 956 282 967 286
rect 907 280 912 281
rect 916 279 937 281
rect 908 275 916 276
rect 920 277 937 279
rect 908 272 920 275
rect 870 261 874 265
rect 831 256 844 260
rect 850 257 874 261
rect 879 262 881 266
rect 761 248 775 252
rect 779 248 780 252
rect 796 252 798 255
rect 831 251 834 256
rect 850 255 854 257
rect 820 247 834 251
rect 837 248 838 252
rect 842 248 843 252
rect 879 253 883 262
rect 908 260 912 272
rect 933 270 937 277
rect 941 275 942 279
rect 946 278 947 279
rect 946 275 958 278
rect 941 274 958 275
rect 954 271 958 274
rect 963 277 967 282
rect 977 279 981 286
rect 977 278 982 279
rect 963 273 970 277
rect 977 274 978 278
rect 985 278 989 299
rect 992 293 1005 294
rect 992 289 995 293
rect 999 289 1001 293
rect 992 288 1005 289
rect 992 281 998 288
rect 1008 282 1012 299
rect 985 274 988 278
rect 992 274 993 278
rect 997 274 998 278
rect 1002 274 1003 278
rect 1008 277 1012 278
rect 977 273 982 274
rect 954 270 959 271
rect 922 264 928 269
rect 933 266 945 270
rect 949 266 950 270
rect 954 266 955 270
rect 922 262 924 264
rect 915 260 924 262
rect 954 265 959 266
rect 954 261 958 265
rect 915 256 928 260
rect 934 257 958 261
rect 908 255 912 256
rect 934 255 938 257
rect 850 250 854 251
rect 859 249 860 253
rect 864 249 883 253
rect 820 243 824 247
rect 837 243 843 248
rect 921 248 922 252
rect 926 248 927 252
rect 963 253 967 273
rect 977 265 981 273
rect 997 269 1003 274
rect 984 265 985 269
rect 989 265 1003 269
rect 1009 268 1013 270
rect 934 250 938 251
rect 943 249 944 253
rect 948 249 967 253
rect 971 262 981 265
rect 971 250 974 262
rect 921 243 927 248
rect 977 256 981 262
rect 977 255 982 256
rect 977 251 978 255
rect 982 251 989 254
rect 977 248 989 251
rect 993 252 997 265
rect 1009 261 1013 264
rect 1000 257 1004 261
rect 1008 257 1013 261
rect 1000 256 1013 257
rect 993 248 1007 252
rect 1011 248 1012 252
rect 744 240 747 243
rect 743 239 747 240
rect 751 239 757 243
rect 761 239 825 243
rect 829 239 878 243
rect 882 239 909 243
rect 913 239 962 243
rect 966 239 979 243
rect 983 239 989 243
rect 993 239 1017 243
rect 743 237 1017 239
rect 724 236 1017 237
rect 727 235 1017 236
rect 727 234 746 235
rect 834 233 878 235
rect 834 229 840 233
rect 844 229 868 233
rect 872 229 878 233
rect 781 227 785 228
rect 725 209 754 214
rect 710 168 715 188
rect 781 186 785 223
rect 838 221 844 229
rect 838 217 839 221
rect 843 217 844 221
rect 849 221 853 222
rect 858 221 864 229
rect 858 217 859 221
rect 863 217 864 221
rect 869 221 874 224
rect 873 217 874 221
rect 849 214 853 217
rect 869 216 874 217
rect 849 210 866 214
rect 797 182 800 201
rect 838 198 842 208
rect 846 203 851 207
rect 862 206 866 210
rect 870 211 886 216
rect 870 206 874 211
rect 846 195 852 199
rect 856 195 859 199
rect 846 189 850 195
rect 862 191 866 202
rect 869 201 883 206
rect 833 186 850 189
rect 854 187 866 191
rect 854 183 858 187
rect 870 186 874 201
rect 869 185 874 186
rect 838 179 839 183
rect 843 179 858 183
rect 861 181 869 183
rect 873 181 874 185
rect 861 179 874 181
rect 954 176 958 183
rect 856 173 857 176
rect 834 172 857 173
rect 861 173 862 176
rect 861 172 868 173
rect 834 169 868 172
rect 872 169 878 173
rect 834 168 878 169
rect 950 168 959 176
rect 710 165 878 168
rect 1040 166 1044 314
rect 1054 311 1407 314
rect 1055 172 1058 311
rect 1233 308 1238 311
rect 1339 308 1343 311
rect 1165 305 1411 308
rect 1165 300 1168 305
rect 1211 299 1214 305
rect 1265 299 1268 305
rect 1321 299 1324 305
rect 1199 288 1202 296
rect 1199 284 1200 288
rect 1182 275 1185 278
rect 1199 262 1202 284
rect 1245 282 1248 295
rect 1245 279 1255 282
rect 1287 279 1290 283
rect 1299 285 1302 295
rect 1299 282 1318 285
rect 1347 285 1350 286
rect 1214 275 1216 278
rect 1236 275 1237 278
rect 1245 270 1248 279
rect 1212 267 1248 270
rect 1212 262 1215 267
rect 1245 262 1248 267
rect 1252 270 1255 279
rect 1266 275 1270 277
rect 1287 276 1291 279
rect 1266 274 1273 275
rect 1299 270 1302 282
rect 1349 281 1350 285
rect 1347 279 1350 281
rect 1323 275 1326 278
rect 1355 275 1358 295
rect 1355 270 1358 271
rect 1266 267 1302 270
rect 1266 262 1269 267
rect 1299 262 1302 267
rect 1322 267 1358 270
rect 1322 262 1325 267
rect 1355 262 1358 267
rect 1165 241 1168 258
rect 1228 241 1231 258
rect 1238 241 1241 244
rect 1282 241 1285 258
rect 1292 241 1295 244
rect 1338 241 1341 258
rect 1366 249 1369 298
rect 1375 299 1378 305
rect 1381 288 1382 292
rect 1379 279 1382 288
rect 1409 284 1412 295
rect 1379 276 1380 279
rect 1398 275 1401 277
rect 1398 274 1404 275
rect 1409 270 1412 280
rect 1376 267 1412 270
rect 1376 262 1379 267
rect 1409 262 1412 267
rect 1423 283 1428 380
rect 1478 366 1484 603
rect 1541 580 1545 699
rect 1676 697 1700 699
rect 1676 696 1717 697
rect 1564 693 1598 696
rect 1564 686 1568 693
rect 1581 663 1584 685
rect 1595 648 1598 693
rect 1676 692 1696 696
rect 1700 693 1717 696
rect 1721 693 1722 697
rect 1729 694 1731 698
rect 1735 694 1743 698
rect 1738 693 1743 694
rect 1676 682 1700 692
rect 1676 678 1696 682
rect 1676 674 1700 678
rect 1705 686 1706 690
rect 1710 686 1711 690
rect 1742 689 1743 693
rect 1705 684 1711 686
rect 1705 680 1706 684
rect 1710 683 1711 684
rect 1721 687 1734 688
rect 1725 683 1734 687
rect 1738 685 1743 689
rect 1747 696 1751 697
rect 1710 680 1718 683
rect 1721 682 1734 683
rect 1747 682 1751 692
rect 1705 677 1718 680
rect 1730 678 1751 682
rect 1756 678 1764 702
rect 1721 677 1725 678
rect 1676 673 1721 674
rect 1676 670 1725 673
rect 1730 674 1734 678
rect 1760 674 1764 678
rect 1612 667 1620 670
rect 1612 663 1616 667
rect 1612 657 1620 663
rect 1625 668 1638 669
rect 1625 664 1628 668
rect 1632 665 1638 668
rect 1642 668 1663 669
rect 1642 665 1651 668
rect 1632 664 1633 665
rect 1650 664 1651 665
rect 1655 665 1663 668
rect 1676 668 1700 670
rect 1730 669 1734 670
rect 1676 667 1696 668
rect 1655 664 1656 665
rect 1625 657 1631 664
rect 1680 664 1696 667
rect 1745 667 1751 674
rect 1720 666 1721 667
rect 1680 663 1700 664
rect 1642 661 1646 662
rect 1676 661 1700 663
rect 1713 663 1721 666
rect 1725 666 1726 667
rect 1743 666 1744 667
rect 1725 663 1744 666
rect 1748 663 1751 667
rect 1713 662 1751 663
rect 1756 668 1764 674
rect 1760 664 1764 668
rect 1612 653 1616 657
rect 1642 653 1646 657
rect 1651 658 1700 661
rect 1734 659 1737 662
rect 1655 657 1700 658
rect 1651 653 1655 654
rect 1612 589 1620 653
rect 1625 649 1646 653
rect 1658 651 1671 654
rect 1625 639 1629 649
rect 1642 648 1655 649
rect 1658 648 1666 651
rect 1625 634 1629 635
rect 1633 642 1638 646
rect 1642 644 1651 648
rect 1642 643 1655 644
rect 1665 647 1666 648
rect 1670 647 1671 651
rect 1665 645 1671 647
rect 1633 638 1634 642
rect 1665 641 1666 645
rect 1670 641 1671 645
rect 1676 653 1700 657
rect 1734 656 1749 659
rect 1680 649 1700 653
rect 1722 652 1725 655
rect 1676 639 1700 649
rect 1633 637 1638 638
rect 1633 633 1640 637
rect 1644 633 1647 637
rect 1654 634 1655 638
rect 1659 635 1676 638
rect 1680 635 1700 639
rect 1659 634 1700 635
rect 1676 631 1700 634
rect 1676 627 1696 631
rect 1628 624 1649 627
rect 1676 615 1700 627
rect 1705 651 1709 652
rect 1705 629 1709 647
rect 1713 648 1750 652
rect 1713 641 1717 648
rect 1728 643 1729 644
rect 1713 636 1717 637
rect 1721 640 1729 643
rect 1733 643 1734 644
rect 1733 640 1742 643
rect 1721 639 1742 640
rect 1721 632 1725 639
rect 1720 631 1725 632
rect 1705 625 1714 629
rect 1724 627 1725 631
rect 1720 626 1725 627
rect 1729 634 1733 635
rect 1710 622 1714 625
rect 1729 622 1733 630
rect 1710 618 1733 622
rect 1738 623 1742 639
rect 1746 633 1750 648
rect 1746 628 1750 629
rect 1756 651 1764 664
rect 1760 647 1764 651
rect 1738 619 1744 623
rect 1748 619 1749 623
rect 1631 612 1652 615
rect 1676 611 1699 615
rect 1703 611 1706 615
rect 1710 611 1711 615
rect 1644 596 1661 599
rect 1658 591 1661 596
rect 1657 590 1671 591
rect 1612 585 1616 589
rect 1632 586 1633 590
rect 1637 586 1653 590
rect 1657 586 1658 590
rect 1662 586 1671 590
rect 1542 558 1550 580
rect 1556 575 1560 576
rect 1556 560 1560 571
rect 1563 568 1566 581
rect 1612 580 1620 585
rect 1606 577 1620 580
rect 1606 576 1629 577
rect 1575 572 1585 576
rect 1594 575 1625 576
rect 1598 574 1625 575
rect 1598 571 1606 574
rect 1594 570 1606 571
rect 1610 572 1625 574
rect 1610 571 1629 572
rect 1633 576 1639 583
rect 1649 582 1653 586
rect 1649 578 1652 582
rect 1656 578 1658 582
rect 1665 579 1671 586
rect 1633 574 1646 576
rect 1610 570 1620 571
rect 1633 570 1637 574
rect 1641 570 1646 574
rect 1563 564 1576 568
rect 1572 562 1576 564
rect 1580 563 1584 568
rect 1542 557 1553 558
rect 1542 553 1549 557
rect 1556 556 1568 560
rect 1542 552 1553 553
rect 1542 546 1550 552
rect 1542 542 1546 546
rect 1542 536 1550 542
rect 1556 545 1560 553
rect 1564 552 1568 556
rect 1587 561 1594 565
rect 1598 561 1599 565
rect 1572 555 1576 558
rect 1587 552 1591 561
rect 1606 556 1620 570
rect 1654 565 1658 578
rect 1676 572 1700 611
rect 1718 605 1722 618
rect 1730 609 1735 613
rect 1739 609 1743 613
rect 1756 612 1764 647
rect 1730 607 1743 609
rect 1705 601 1711 604
rect 1718 601 1720 605
rect 1724 601 1727 605
rect 1705 597 1706 601
rect 1710 597 1711 601
rect 1723 597 1727 601
rect 1737 600 1743 607
rect 1747 611 1764 612
rect 1751 607 1764 611
rect 1747 606 1764 607
rect 1756 598 1764 606
rect 1705 593 1714 597
rect 1718 593 1719 597
rect 1723 593 1739 597
rect 1743 593 1744 597
rect 1760 594 1764 598
rect 1705 592 1719 593
rect 1709 578 1748 581
rect 1752 578 1753 581
rect 1665 568 1666 572
rect 1670 568 1673 572
rect 1677 568 1700 572
rect 1627 560 1628 564
rect 1632 560 1638 564
rect 1564 548 1579 552
rect 1583 548 1591 552
rect 1594 555 1620 556
rect 1598 551 1620 555
rect 1594 550 1620 551
rect 1606 546 1620 550
rect 1556 541 1558 545
rect 1562 544 1563 545
rect 1593 544 1594 545
rect 1562 541 1580 544
rect 1556 540 1580 541
rect 1584 541 1594 544
rect 1598 541 1601 545
rect 1584 540 1601 541
rect 1610 542 1620 546
rect 1606 536 1620 542
rect 1612 532 1616 536
rect 1612 505 1620 532
rect 1626 554 1630 555
rect 1626 535 1630 550
rect 1634 544 1638 560
rect 1643 561 1666 565
rect 1643 553 1647 561
rect 1662 558 1666 561
rect 1643 548 1647 549
rect 1651 556 1656 557
rect 1651 552 1652 556
rect 1662 554 1671 558
rect 1651 551 1656 552
rect 1651 544 1655 551
rect 1634 543 1655 544
rect 1634 540 1643 543
rect 1642 539 1643 540
rect 1647 540 1655 543
rect 1659 546 1663 547
rect 1647 539 1648 540
rect 1659 535 1663 542
rect 1626 533 1663 535
rect 1626 531 1639 533
rect 1643 531 1663 533
rect 1667 536 1671 554
rect 1667 531 1671 532
rect 1676 556 1700 568
rect 1680 552 1700 556
rect 1676 547 1700 552
rect 1676 543 1696 547
rect 1676 531 1700 543
rect 1705 567 1709 568
rect 1705 545 1709 563
rect 1713 566 1733 568
rect 1737 566 1750 568
rect 1713 564 1750 566
rect 1713 557 1717 564
rect 1728 559 1729 560
rect 1713 552 1717 553
rect 1721 556 1729 559
rect 1733 559 1734 560
rect 1733 556 1742 559
rect 1721 555 1742 556
rect 1721 548 1725 555
rect 1720 547 1725 548
rect 1705 541 1714 545
rect 1724 543 1725 547
rect 1720 542 1725 543
rect 1729 550 1733 551
rect 1710 538 1714 541
rect 1729 538 1733 546
rect 1710 534 1733 538
rect 1738 539 1742 555
rect 1746 549 1750 564
rect 1746 544 1750 545
rect 1756 567 1764 594
rect 1774 578 1790 581
rect 1760 563 1764 567
rect 1756 557 1770 563
rect 1787 559 1790 578
rect 1828 563 1834 755
rect 1756 553 1766 557
rect 1775 558 1820 559
rect 1775 554 1778 558
rect 1782 555 1814 558
rect 1782 554 1783 555
rect 1813 554 1814 555
rect 1818 554 1820 558
rect 1756 549 1770 553
rect 1756 548 1782 549
rect 1756 544 1778 548
rect 1756 543 1782 544
rect 1785 547 1793 551
rect 1797 547 1812 551
rect 1738 535 1744 539
rect 1748 535 1749 539
rect 1676 527 1699 531
rect 1703 527 1706 531
rect 1710 527 1711 531
rect 1625 520 1652 521
rect 1628 517 1648 520
rect 1657 506 1671 507
rect 1612 501 1616 505
rect 1632 502 1633 506
rect 1637 502 1653 506
rect 1657 502 1658 506
rect 1662 502 1671 506
rect 1612 493 1620 501
rect 1612 492 1629 493
rect 1612 488 1625 492
rect 1612 487 1629 488
rect 1633 492 1639 499
rect 1649 498 1653 502
rect 1665 498 1666 502
rect 1670 498 1671 502
rect 1649 494 1652 498
rect 1656 494 1658 498
rect 1665 495 1671 498
rect 1633 490 1646 492
rect 1495 468 1566 472
rect 1496 438 1531 442
rect 1478 361 1502 366
rect 1433 348 1483 352
rect 1433 298 1437 348
rect 1447 344 1453 348
rect 1457 344 1483 348
rect 1462 339 1468 344
rect 1462 335 1463 339
rect 1467 335 1468 339
rect 1474 338 1479 339
rect 1478 334 1479 338
rect 1474 331 1479 334
rect 1451 327 1452 331
rect 1456 327 1471 331
rect 1451 322 1463 323
rect 1451 318 1455 322
rect 1459 318 1463 322
rect 1451 317 1463 318
rect 1467 322 1471 327
rect 1478 327 1479 331
rect 1474 326 1479 327
rect 1448 314 1455 317
rect 1451 309 1455 314
rect 1467 306 1471 318
rect 1475 315 1479 326
rect 1475 312 1489 315
rect 1475 306 1479 312
rect 1451 302 1452 306
rect 1456 302 1471 306
rect 1474 305 1479 306
rect 1478 301 1479 305
rect 1474 298 1479 301
rect 1433 295 1435 298
rect 1466 294 1474 298
rect 1478 294 1479 298
rect 1466 293 1479 294
rect 1447 284 1453 288
rect 1457 284 1463 288
rect 1467 284 1483 288
rect 1447 283 1483 284
rect 1423 280 1483 283
rect 1348 241 1351 244
rect 1392 241 1395 258
rect 1402 241 1405 244
rect 1423 241 1428 280
rect 1475 263 1478 280
rect 1474 259 1478 263
rect 1449 255 1485 259
rect 1449 251 1455 255
rect 1459 251 1465 255
rect 1469 251 1485 255
rect 1468 245 1481 246
rect 1468 241 1476 245
rect 1480 241 1481 245
rect 1063 238 1429 241
rect 1079 219 1082 238
rect 1162 236 1429 238
rect 1476 238 1481 241
rect 1124 221 1128 223
rect 1162 219 1165 236
rect 1174 229 1205 232
rect 1124 204 1128 215
rect 1107 200 1110 203
rect 1124 194 1127 204
rect 1179 199 1182 202
rect 1124 190 1125 194
rect 1196 193 1199 215
rect 1202 203 1205 229
rect 1225 219 1228 236
rect 1235 233 1238 236
rect 1279 219 1282 236
rect 1289 233 1292 236
rect 1335 219 1338 236
rect 1345 233 1348 236
rect 1389 219 1392 236
rect 1399 233 1402 236
rect 1209 210 1212 215
rect 1242 210 1245 215
rect 1209 207 1245 210
rect 1202 200 1207 203
rect 1211 199 1213 202
rect 1233 199 1234 202
rect 1242 198 1245 207
rect 1263 210 1266 215
rect 1296 210 1299 215
rect 1263 207 1299 210
rect 1319 210 1322 215
rect 1352 210 1355 215
rect 1319 207 1355 210
rect 1249 198 1252 207
rect 1263 202 1270 203
rect 1263 200 1267 202
rect 1284 198 1288 201
rect 1242 195 1252 198
rect 1124 182 1127 190
rect 1196 189 1197 193
rect 1196 181 1199 189
rect 1242 182 1245 195
rect 1284 194 1287 198
rect 1296 195 1299 207
rect 1352 206 1355 207
rect 1362 214 1364 218
rect 1320 199 1323 202
rect 1296 192 1315 195
rect 1296 182 1299 192
rect 1344 196 1347 198
rect 1332 188 1335 194
rect 1346 192 1347 196
rect 1344 191 1347 192
rect 1309 185 1335 188
rect 1352 182 1355 202
rect 1090 172 1093 178
rect 1362 179 1366 214
rect 1373 210 1376 215
rect 1406 210 1409 215
rect 1373 207 1409 210
rect 1376 198 1377 201
rect 1395 202 1401 203
rect 1395 200 1398 202
rect 1376 189 1379 198
rect 1406 197 1409 207
rect 1378 185 1379 189
rect 1406 182 1409 193
rect 1162 172 1165 177
rect 1208 172 1211 178
rect 1262 172 1265 178
rect 1318 172 1321 178
rect 1365 177 1366 179
rect 1372 172 1375 178
rect 1055 169 1409 172
rect 1234 166 1239 169
rect 1340 166 1344 169
rect 710 164 834 165
rect 1040 162 1102 166
rect 771 153 1086 158
rect 393 138 399 146
rect 393 134 394 138
rect 398 134 399 138
rect 404 140 408 141
rect 413 140 419 146
rect 454 140 465 143
rect 413 136 414 140
rect 418 136 419 140
rect 383 133 388 134
rect 383 129 384 133
rect 404 133 408 136
rect 383 126 388 129
rect 383 122 384 126
rect 383 121 388 122
rect 391 129 404 131
rect 391 127 408 129
rect 415 129 446 133
rect 383 120 387 121
rect 347 116 387 120
rect 344 104 374 107
rect 383 103 387 116
rect 391 116 395 127
rect 406 120 411 124
rect 415 120 419 129
rect 398 112 401 116
rect 405 112 412 116
rect 391 108 395 112
rect 391 104 403 108
rect 407 107 412 112
rect 383 102 388 103
rect 383 98 384 102
rect 388 98 395 101
rect 383 95 395 98
rect 399 100 403 104
rect 406 103 422 107
rect 399 96 414 100
rect 418 96 419 100
rect 442 96 446 129
rect 462 130 465 140
rect 486 138 492 146
rect 486 134 487 138
rect 491 134 492 138
rect 497 140 501 141
rect 506 140 512 146
rect 506 136 507 140
rect 511 136 512 140
rect 573 138 579 146
rect 552 137 568 138
rect 476 133 481 134
rect 476 130 477 133
rect 462 129 477 130
rect 497 133 501 136
rect 462 127 481 129
rect 476 126 481 127
rect 476 122 477 126
rect 476 121 481 122
rect 484 129 497 131
rect 484 127 501 129
rect 476 103 480 121
rect 484 116 488 127
rect 508 124 512 133
rect 556 133 568 137
rect 573 134 574 138
rect 578 134 579 138
rect 584 140 588 141
rect 593 140 599 146
rect 699 143 1074 146
rect 824 142 1074 143
rect 593 136 594 140
rect 598 136 599 140
rect 556 132 564 133
rect 563 129 564 132
rect 584 133 588 136
rect 563 126 568 129
rect 499 120 504 124
rect 508 120 519 124
rect 563 122 564 126
rect 563 121 568 122
rect 571 129 584 131
rect 571 127 588 129
rect 491 112 494 116
rect 498 112 505 116
rect 484 108 488 112
rect 484 104 496 108
rect 476 102 481 103
rect 476 98 477 102
rect 481 98 488 101
rect 476 95 488 98
rect 492 100 496 104
rect 500 107 505 112
rect 500 103 515 107
rect 563 103 567 121
rect 571 116 575 127
rect 595 124 599 133
rect 1045 131 1048 133
rect 1045 128 1052 131
rect 586 120 591 124
rect 595 120 608 124
rect 578 112 581 116
rect 585 112 592 116
rect 571 108 575 112
rect 571 104 583 108
rect 563 102 568 103
rect 492 96 507 100
rect 511 96 512 100
rect 563 98 564 102
rect 568 98 575 101
rect 563 95 575 98
rect 579 100 583 104
rect 587 106 592 112
rect 1045 108 1048 128
rect 587 103 600 106
rect 1026 107 1049 108
rect 605 103 1049 107
rect 579 96 594 100
rect 598 96 599 100
rect 379 86 385 90
rect 389 86 395 90
rect 399 86 423 90
rect 472 86 478 90
rect 482 86 488 90
rect 492 86 516 90
rect 373 85 516 86
rect 559 86 565 90
rect 569 86 575 90
rect 579 86 603 90
rect 559 85 603 86
rect 373 83 603 85
rect 379 82 423 83
rect 472 82 603 83
rect 1068 71 1073 142
rect 1083 84 1086 153
rect 1098 95 1102 162
rect 1166 163 1412 166
rect 1166 158 1169 163
rect 1114 153 1148 157
rect 1212 157 1215 163
rect 1266 157 1269 163
rect 1322 157 1325 163
rect 1200 146 1203 154
rect 1200 142 1201 146
rect 1183 133 1186 136
rect 1200 120 1203 142
rect 1246 140 1249 153
rect 1246 137 1256 140
rect 1288 137 1291 141
rect 1300 143 1303 153
rect 1300 140 1319 143
rect 1348 143 1351 144
rect 1215 133 1217 136
rect 1237 133 1238 136
rect 1246 128 1249 137
rect 1213 125 1249 128
rect 1213 120 1216 125
rect 1246 120 1249 125
rect 1253 128 1256 137
rect 1267 133 1271 135
rect 1288 134 1292 137
rect 1267 132 1274 133
rect 1300 128 1303 140
rect 1350 139 1351 143
rect 1348 137 1351 139
rect 1324 133 1327 136
rect 1356 133 1359 153
rect 1356 128 1359 129
rect 1267 125 1303 128
rect 1267 120 1270 125
rect 1300 120 1303 125
rect 1323 125 1359 128
rect 1323 120 1326 125
rect 1356 120 1359 125
rect 1166 97 1169 116
rect 1229 97 1232 116
rect 1239 97 1242 102
rect 1283 97 1286 116
rect 1293 97 1296 102
rect 1339 97 1342 116
rect 1365 105 1368 156
rect 1376 157 1379 163
rect 1382 146 1383 150
rect 1380 137 1383 146
rect 1410 142 1413 153
rect 1380 134 1381 137
rect 1399 133 1402 135
rect 1399 132 1405 133
rect 1410 128 1413 138
rect 1377 125 1413 128
rect 1377 120 1380 125
rect 1410 120 1413 125
rect 1349 97 1352 102
rect 1393 97 1396 116
rect 1424 105 1429 236
rect 1453 233 1454 237
rect 1458 233 1473 237
rect 1480 234 1481 238
rect 1476 233 1481 234
rect 1447 228 1458 230
rect 1451 224 1458 228
rect 1453 222 1458 224
rect 1453 221 1465 222
rect 1453 217 1457 221
rect 1461 217 1465 221
rect 1453 216 1465 217
rect 1469 221 1473 233
rect 1469 212 1473 217
rect 1477 224 1481 233
rect 1497 229 1502 361
rect 1560 354 1564 468
rect 1590 332 1593 457
rect 1514 328 1593 332
rect 1612 452 1620 487
rect 1633 486 1637 490
rect 1641 486 1646 490
rect 1654 481 1658 494
rect 1676 488 1700 527
rect 1718 521 1722 534
rect 1756 529 1770 543
rect 1785 538 1789 547
rect 1800 541 1804 544
rect 1777 534 1778 538
rect 1782 534 1789 538
rect 1808 543 1812 547
rect 1816 546 1820 554
rect 1826 557 1834 563
rect 1830 553 1834 557
rect 1826 547 1834 553
rect 1823 546 1834 547
rect 1808 539 1820 543
rect 1827 542 1834 546
rect 1823 541 1834 542
rect 1792 531 1796 536
rect 1800 535 1804 537
rect 1800 531 1813 535
rect 1730 525 1735 529
rect 1739 525 1743 529
rect 1756 528 1766 529
rect 1730 523 1743 525
rect 1705 513 1711 520
rect 1718 517 1720 521
rect 1724 517 1727 521
rect 1723 513 1727 517
rect 1737 516 1743 523
rect 1747 527 1766 528
rect 1751 525 1766 527
rect 1770 528 1782 529
rect 1770 525 1778 528
rect 1751 524 1778 525
rect 1751 523 1782 524
rect 1791 523 1801 527
rect 1747 522 1770 523
rect 1756 519 1770 522
rect 1756 514 1764 519
rect 1810 518 1813 531
rect 1816 528 1820 539
rect 1816 523 1820 524
rect 1826 519 1834 541
rect 1705 509 1714 513
rect 1718 509 1719 513
rect 1723 509 1739 513
rect 1743 509 1744 513
rect 1760 510 1764 514
rect 1705 508 1719 509
rect 1715 503 1718 508
rect 1756 505 1764 510
rect 1715 500 1732 503
rect 1756 502 1778 505
rect 1665 484 1666 488
rect 1670 484 1673 488
rect 1677 484 1700 488
rect 1627 476 1628 480
rect 1632 476 1638 480
rect 1600 335 1603 450
rect 1612 448 1616 452
rect 1612 435 1620 448
rect 1626 470 1630 471
rect 1626 451 1630 466
rect 1634 460 1638 476
rect 1643 477 1666 481
rect 1643 469 1647 477
rect 1662 474 1666 477
rect 1643 464 1647 465
rect 1651 472 1656 473
rect 1651 468 1652 472
rect 1662 470 1671 474
rect 1651 467 1656 468
rect 1651 460 1655 467
rect 1634 459 1655 460
rect 1634 456 1643 459
rect 1642 455 1643 456
rect 1647 456 1655 459
rect 1659 462 1663 463
rect 1647 455 1648 456
rect 1659 451 1663 458
rect 1626 447 1663 451
rect 1667 452 1671 470
rect 1667 447 1671 448
rect 1676 472 1700 484
rect 1680 468 1700 472
rect 1676 465 1700 468
rect 1756 493 1770 502
rect 1778 493 1779 500
rect 1756 490 1779 493
rect 1676 464 1717 465
rect 1676 460 1696 464
rect 1700 461 1717 464
rect 1721 461 1722 465
rect 1729 462 1732 466
rect 1736 462 1743 466
rect 1738 461 1743 462
rect 1676 450 1700 460
rect 1649 444 1653 447
rect 1627 440 1642 443
rect 1676 446 1696 450
rect 1676 442 1700 446
rect 1705 454 1706 458
rect 1710 454 1711 458
rect 1742 457 1743 461
rect 1705 452 1711 454
rect 1705 448 1706 452
rect 1710 451 1711 452
rect 1721 455 1734 456
rect 1725 451 1734 455
rect 1738 453 1743 457
rect 1747 464 1751 465
rect 1710 448 1718 451
rect 1721 450 1734 451
rect 1747 450 1751 460
rect 1705 445 1718 448
rect 1730 446 1751 450
rect 1756 446 1770 490
rect 1788 484 1823 485
rect 1788 480 1818 484
rect 1721 445 1725 446
rect 1676 441 1721 442
rect 1639 437 1642 440
rect 1676 438 1725 441
rect 1730 442 1734 446
rect 1760 442 1770 446
rect 1612 431 1616 435
rect 1612 425 1620 431
rect 1625 436 1663 437
rect 1625 432 1628 436
rect 1632 433 1651 436
rect 1632 432 1633 433
rect 1650 432 1651 433
rect 1655 433 1663 436
rect 1676 436 1700 438
rect 1730 437 1734 438
rect 1676 435 1696 436
rect 1655 432 1656 433
rect 1625 425 1631 432
rect 1680 432 1696 435
rect 1745 435 1751 442
rect 1720 434 1721 435
rect 1680 431 1700 432
rect 1642 429 1646 430
rect 1676 429 1700 431
rect 1713 431 1721 434
rect 1725 434 1726 435
rect 1743 434 1744 435
rect 1725 431 1734 434
rect 1713 430 1734 431
rect 1738 431 1744 434
rect 1748 431 1751 435
rect 1738 430 1751 431
rect 1756 437 1770 442
rect 1756 436 1810 437
rect 1760 432 1810 436
rect 1756 429 1770 432
rect 1612 421 1616 425
rect 1642 421 1646 425
rect 1651 426 1700 429
rect 1655 425 1700 426
rect 1651 421 1655 422
rect 1612 397 1620 421
rect 1625 417 1646 421
rect 1658 419 1671 422
rect 1625 407 1629 417
rect 1642 416 1655 417
rect 1658 416 1666 419
rect 1625 402 1629 403
rect 1633 410 1638 414
rect 1642 412 1651 416
rect 1642 411 1655 412
rect 1665 415 1666 416
rect 1670 415 1671 419
rect 1665 413 1671 415
rect 1633 406 1634 410
rect 1665 409 1666 413
rect 1670 409 1671 413
rect 1676 421 1700 425
rect 1680 417 1700 421
rect 1676 407 1700 417
rect 1760 415 1770 429
rect 1760 412 1762 415
rect 1633 405 1638 406
rect 1633 401 1641 405
rect 1645 401 1647 405
rect 1654 402 1655 406
rect 1659 403 1676 406
rect 1680 404 1700 407
rect 1680 403 1684 404
rect 1659 402 1684 403
rect 1676 398 1684 402
rect 1690 400 1700 404
rect 1831 400 1835 519
rect 1690 398 1835 400
rect 1676 397 1835 398
rect 1614 369 1619 397
rect 1692 396 1835 397
rect 1811 395 1835 396
rect 1715 384 1758 389
rect 1809 387 1814 388
rect 1614 368 1740 369
rect 1614 363 1735 368
rect 1684 350 1685 352
rect 1771 354 1772 357
rect 1776 354 1801 357
rect 1684 346 1690 350
rect 1684 341 1692 346
rect 1748 345 1756 346
rect 1809 345 1814 382
rect 1684 340 1709 341
rect 1684 336 1688 340
rect 1692 337 1709 340
rect 1713 337 1714 341
rect 1721 338 1723 342
rect 1727 338 1735 342
rect 1730 337 1735 338
rect 1600 325 1604 335
rect 1684 326 1692 336
rect 1684 322 1688 326
rect 1684 318 1692 322
rect 1697 330 1698 334
rect 1702 330 1703 334
rect 1734 333 1735 337
rect 1697 328 1703 330
rect 1697 324 1698 328
rect 1702 327 1703 328
rect 1713 331 1726 332
rect 1717 327 1726 331
rect 1730 329 1735 333
rect 1739 340 1743 341
rect 1702 324 1710 327
rect 1713 326 1726 327
rect 1739 326 1743 336
rect 1697 321 1710 324
rect 1722 322 1743 326
rect 1748 340 1814 345
rect 1748 322 1756 340
rect 1713 321 1717 322
rect 1684 317 1713 318
rect 1684 314 1717 317
rect 1722 318 1726 322
rect 1752 318 1756 322
rect 1684 312 1692 314
rect 1722 313 1726 314
rect 1684 308 1688 312
rect 1737 311 1743 318
rect 1712 310 1713 311
rect 1510 294 1650 296
rect 1510 292 1645 294
rect 1684 275 1692 308
rect 1705 307 1713 310
rect 1717 310 1718 311
rect 1735 310 1736 311
rect 1717 307 1736 310
rect 1740 307 1743 311
rect 1705 306 1743 307
rect 1748 312 1756 318
rect 1752 308 1756 312
rect 1726 303 1729 306
rect 1726 300 1741 303
rect 1711 296 1714 299
rect 1684 271 1688 275
rect 1684 259 1692 271
rect 1697 295 1701 296
rect 1697 273 1701 291
rect 1705 292 1742 296
rect 1705 285 1709 292
rect 1720 287 1721 288
rect 1705 280 1709 281
rect 1713 284 1721 287
rect 1725 287 1726 288
rect 1725 284 1734 287
rect 1713 283 1734 284
rect 1713 276 1717 283
rect 1712 275 1717 276
rect 1697 269 1706 273
rect 1716 271 1717 275
rect 1712 270 1717 271
rect 1721 278 1725 279
rect 1702 266 1706 269
rect 1721 266 1725 274
rect 1702 262 1725 266
rect 1730 267 1734 283
rect 1738 277 1742 292
rect 1738 272 1742 273
rect 1748 295 1756 308
rect 1752 291 1756 295
rect 1730 263 1736 267
rect 1740 263 1741 267
rect 1684 255 1691 259
rect 1695 255 1698 259
rect 1702 255 1703 259
rect 1477 221 1488 224
rect 1477 213 1481 221
rect 1453 208 1454 212
rect 1458 208 1473 212
rect 1476 212 1481 213
rect 1480 208 1481 212
rect 1476 205 1481 208
rect 1464 200 1465 204
rect 1469 200 1470 204
rect 1480 201 1481 205
rect 1476 200 1481 201
rect 1497 216 1501 229
rect 1646 225 1652 227
rect 1508 224 1652 225
rect 1508 221 1647 224
rect 1646 220 1647 221
rect 1651 220 1652 224
rect 1464 195 1470 200
rect 1449 191 1455 195
rect 1459 191 1485 195
rect 1449 187 1485 191
rect 1478 173 1481 187
rect 1451 169 1487 173
rect 1451 165 1457 169
rect 1461 165 1487 169
rect 1466 160 1472 165
rect 1466 156 1467 160
rect 1471 156 1472 160
rect 1478 159 1483 160
rect 1482 155 1483 159
rect 1478 152 1483 155
rect 1455 148 1456 152
rect 1460 148 1475 152
rect 1455 143 1467 144
rect 1455 142 1459 143
rect 1444 139 1459 142
rect 1463 139 1467 143
rect 1455 138 1467 139
rect 1471 143 1475 148
rect 1482 148 1483 152
rect 1478 147 1483 148
rect 1455 130 1459 138
rect 1471 127 1475 139
rect 1479 139 1483 147
rect 1479 135 1488 139
rect 1492 135 1493 139
rect 1479 127 1483 135
rect 1455 123 1456 127
rect 1460 123 1475 127
rect 1478 126 1483 127
rect 1482 122 1483 126
rect 1478 119 1483 122
rect 1470 115 1478 119
rect 1482 115 1483 119
rect 1470 114 1483 115
rect 1497 112 1502 216
rect 1684 191 1692 255
rect 1710 249 1714 262
rect 1722 253 1727 257
rect 1731 253 1735 257
rect 1748 256 1756 291
rect 1773 276 1777 317
rect 1858 311 1861 1097
rect 1872 1083 1922 1086
rect 1872 783 1877 1083
rect 1905 998 1908 1009
rect 1905 882 1908 989
rect 1929 967 1932 1133
rect 1948 1097 2009 1100
rect 1929 962 1932 963
rect 1999 928 2003 1097
rect 2009 943 2012 1082
rect 2211 1019 2214 1020
rect 2211 1016 3004 1019
rect 2009 940 2088 943
rect 1999 924 2005 928
rect 2083 894 2087 940
rect 2211 892 2214 1016
rect 2289 999 3011 1002
rect 2289 928 2292 999
rect 2635 983 3011 986
rect 2632 939 2635 982
rect 2708 951 2711 962
rect 2800 949 2803 966
rect 2851 936 2975 937
rect 2674 935 2774 936
rect 2807 935 2975 936
rect 2491 934 2620 935
rect 2447 932 2620 934
rect 2641 933 2975 935
rect 2641 932 2851 933
rect 2447 931 2813 932
rect 2447 930 2491 931
rect 2447 926 2453 930
rect 2457 927 2491 930
rect 2457 926 2464 927
rect 2463 923 2464 926
rect 2468 926 2491 927
rect 2610 929 2813 931
rect 2468 923 2469 926
rect 2451 918 2464 920
rect 2451 914 2452 918
rect 2456 916 2464 918
rect 2467 916 2482 920
rect 2486 916 2487 920
rect 2451 913 2456 914
rect 2451 896 2455 913
rect 2467 912 2471 916
rect 2451 883 2455 892
rect 2459 908 2471 912
rect 2475 910 2492 913
rect 2459 897 2463 908
rect 2475 904 2479 910
rect 2610 911 2615 929
rect 2674 928 2690 929
rect 2689 925 2690 928
rect 2694 928 2725 929
rect 2694 925 2695 928
rect 2724 925 2725 928
rect 2729 928 2747 929
rect 2729 925 2730 928
rect 2724 922 2730 925
rect 2746 925 2747 928
rect 2751 928 2774 929
rect 2807 928 2813 929
rect 2817 929 2851 932
rect 2817 928 2824 929
rect 2751 925 2752 928
rect 2823 925 2824 928
rect 2828 928 2851 929
rect 2828 925 2829 928
rect 2746 922 2752 925
rect 2678 918 2691 922
rect 2724 918 2725 922
rect 2729 918 2730 922
rect 2737 921 2741 922
rect 2678 917 2683 918
rect 2678 913 2679 917
rect 2694 914 2718 918
rect 2746 918 2747 922
rect 2751 918 2752 922
rect 2811 920 2824 922
rect 2737 914 2741 917
rect 2757 914 2763 915
rect 2466 900 2469 904
rect 2473 900 2479 904
rect 2459 889 2463 893
rect 2474 892 2479 896
rect 2483 891 2487 901
rect 2574 892 2596 895
rect 2459 885 2476 889
rect 1905 879 2379 882
rect 2451 882 2456 883
rect 2472 882 2476 885
rect 2451 878 2452 882
rect 2451 875 2456 878
rect 2461 878 2462 882
rect 2466 878 2467 882
rect 1926 870 2380 873
rect 1922 868 1968 870
rect 2461 870 2467 878
rect 2472 877 2476 878
rect 2481 878 2482 882
rect 2486 878 2487 882
rect 2481 870 2487 878
rect 1872 782 1878 783
rect 1822 308 1862 311
rect 1784 291 1837 292
rect 1873 291 1878 782
rect 1886 775 1891 776
rect 1886 769 1905 775
rect 1886 715 1891 769
rect 1886 493 1892 715
rect 1922 644 1930 868
rect 2447 866 2453 870
rect 2457 866 2481 870
rect 2485 866 2491 870
rect 2447 864 2491 866
rect 2308 862 2581 864
rect 2274 860 2581 862
rect 2274 857 2332 860
rect 1972 848 2005 852
rect 2010 848 2011 852
rect 1972 847 2011 848
rect 1972 804 1975 847
rect 1940 800 1975 804
rect 1940 799 1973 800
rect 2132 799 2135 819
rect 2211 799 2214 848
rect 1940 772 1944 799
rect 1951 791 2263 792
rect 1951 789 2261 791
rect 1951 788 2206 789
rect 1951 784 1987 788
rect 1991 784 2001 788
rect 2005 784 2015 788
rect 2019 785 2098 788
rect 2019 784 2082 785
rect 1951 673 1955 784
rect 1963 747 1967 776
rect 1966 743 1967 747
rect 1985 764 1989 771
rect 1985 763 1990 764
rect 1985 759 1986 763
rect 1993 763 1997 784
rect 2000 778 2013 779
rect 2000 774 2003 778
rect 2007 774 2009 778
rect 2000 773 2013 774
rect 2000 766 2006 773
rect 2016 767 2020 784
rect 2086 784 2098 785
rect 2102 785 2182 788
rect 2102 784 2166 785
rect 2063 773 2075 779
rect 2082 778 2086 781
rect 2170 784 2182 785
rect 2186 784 2206 788
rect 2217 788 2261 789
rect 2096 775 2118 779
rect 2122 775 2123 779
rect 2147 778 2159 779
rect 2132 775 2152 778
rect 2096 774 2100 775
rect 2082 773 2086 774
rect 2063 770 2068 773
rect 1993 759 1996 763
rect 2000 759 2001 763
rect 2005 759 2006 763
rect 2010 759 2011 763
rect 2016 762 2020 763
rect 2063 769 2064 770
rect 2059 766 2064 769
rect 2089 770 2100 774
rect 2089 766 2093 770
rect 2107 767 2108 771
rect 2112 767 2123 771
rect 1985 758 1990 759
rect 1985 750 1989 758
rect 2005 754 2011 759
rect 1992 750 1993 754
rect 1997 750 2011 754
rect 2017 752 2021 755
rect 2055 752 2058 766
rect 2063 765 2068 766
rect 2072 764 2093 766
rect 1985 741 1989 746
rect 1985 740 1990 741
rect 1985 736 1986 740
rect 1990 736 1997 739
rect 1985 733 1997 736
rect 2001 737 2005 750
rect 2064 760 2072 761
rect 2076 762 2093 764
rect 2064 757 2076 760
rect 2017 746 2021 748
rect 2008 742 2012 746
rect 2016 742 2021 746
rect 2008 741 2021 742
rect 2064 745 2068 757
rect 2089 755 2093 762
rect 2097 760 2098 764
rect 2102 763 2103 764
rect 2102 760 2114 763
rect 2097 759 2114 760
rect 2110 756 2114 759
rect 2110 755 2115 756
rect 2078 749 2084 754
rect 2089 751 2101 755
rect 2105 751 2106 755
rect 2110 751 2111 755
rect 2078 747 2080 749
rect 2071 745 2080 747
rect 2110 750 2115 751
rect 2119 751 2123 767
rect 2110 746 2114 750
rect 2071 741 2084 745
rect 2090 742 2114 746
rect 2119 747 2121 751
rect 2064 740 2068 741
rect 2090 740 2094 742
rect 2001 733 2015 737
rect 2019 733 2020 737
rect 2077 733 2078 737
rect 2082 733 2083 737
rect 2119 738 2123 747
rect 2090 735 2094 736
rect 2099 734 2100 738
rect 2104 734 2123 738
rect 2132 735 2135 775
rect 2147 774 2152 775
rect 2156 774 2159 778
rect 2147 773 2159 774
rect 2166 778 2170 781
rect 2217 784 2219 788
rect 2223 784 2233 788
rect 2237 784 2247 788
rect 2251 786 2261 788
rect 2251 784 2257 786
rect 2180 775 2202 779
rect 2206 775 2207 779
rect 2180 774 2184 775
rect 2166 773 2170 774
rect 2147 770 2152 773
rect 2147 766 2148 770
rect 2173 770 2184 774
rect 2173 766 2177 770
rect 2191 767 2192 771
rect 2196 767 2207 771
rect 2147 765 2152 766
rect 2156 764 2177 766
rect 2148 760 2156 761
rect 2160 762 2177 764
rect 2148 757 2160 760
rect 2148 745 2152 757
rect 2173 755 2177 762
rect 2181 760 2182 764
rect 2186 763 2187 764
rect 2186 760 2198 763
rect 2181 759 2198 760
rect 2194 756 2198 759
rect 2203 759 2207 767
rect 2210 759 2213 782
rect 2203 756 2213 759
rect 2217 764 2221 771
rect 2217 763 2222 764
rect 2217 759 2218 763
rect 2225 763 2229 784
rect 2232 778 2245 779
rect 2232 774 2235 778
rect 2239 774 2241 778
rect 2232 773 2245 774
rect 2232 766 2238 773
rect 2248 767 2252 784
rect 2225 759 2228 763
rect 2232 759 2233 763
rect 2237 759 2238 763
rect 2242 759 2243 763
rect 2248 762 2252 763
rect 2217 758 2222 759
rect 2194 755 2199 756
rect 2162 749 2168 754
rect 2173 751 2185 755
rect 2189 751 2190 755
rect 2194 751 2195 755
rect 2162 747 2164 749
rect 2155 745 2164 747
rect 2194 750 2199 751
rect 2194 746 2198 750
rect 2155 741 2168 745
rect 2174 742 2198 746
rect 2148 740 2152 741
rect 2174 740 2178 742
rect 2077 728 2083 733
rect 2161 733 2162 737
rect 2166 733 2167 737
rect 2203 738 2207 756
rect 2217 750 2221 758
rect 2237 754 2243 759
rect 2224 750 2225 754
rect 2229 750 2243 754
rect 2249 753 2253 755
rect 2174 735 2178 736
rect 2183 734 2184 738
rect 2188 734 2207 738
rect 2211 747 2221 750
rect 2211 735 2214 747
rect 2161 728 2167 733
rect 2217 741 2221 747
rect 2217 740 2222 741
rect 2217 736 2218 740
rect 2222 736 2229 739
rect 2217 733 2229 736
rect 2233 737 2237 750
rect 2249 746 2253 749
rect 2240 742 2244 746
rect 2248 742 2253 746
rect 2240 741 2253 742
rect 2274 741 2280 857
rect 2308 856 2332 857
rect 2336 856 2342 860
rect 2346 856 2359 860
rect 2363 856 2412 860
rect 2416 856 2443 860
rect 2447 856 2496 860
rect 2500 856 2564 860
rect 2568 856 2574 860
rect 2578 856 2581 860
rect 2313 847 2314 851
rect 2318 847 2332 851
rect 2312 842 2325 843
rect 2312 838 2317 842
rect 2321 838 2325 842
rect 2312 835 2316 838
rect 2328 834 2332 847
rect 2336 848 2348 851
rect 2336 845 2343 848
rect 2347 844 2348 848
rect 2343 843 2348 844
rect 2344 837 2348 843
rect 2398 851 2404 856
rect 2351 837 2354 849
rect 2344 834 2354 837
rect 2358 846 2377 850
rect 2381 846 2382 850
rect 2387 848 2391 849
rect 2312 829 2316 831
rect 2322 830 2336 834
rect 2340 830 2341 834
rect 2322 825 2328 830
rect 2344 826 2348 834
rect 2343 825 2348 826
rect 2313 821 2317 822
rect 2322 821 2323 825
rect 2327 821 2328 825
rect 2332 821 2333 825
rect 2337 821 2340 825
rect 2313 800 2317 817
rect 2327 811 2333 818
rect 2320 810 2333 811
rect 2324 806 2326 810
rect 2330 806 2333 810
rect 2320 805 2333 806
rect 2336 800 2340 821
rect 2347 821 2348 825
rect 2343 820 2348 821
rect 2344 813 2348 820
rect 2358 817 2362 846
rect 2398 847 2399 851
rect 2403 847 2404 851
rect 2482 851 2488 856
rect 2442 846 2461 850
rect 2465 846 2466 850
rect 2471 848 2475 849
rect 2387 842 2391 844
rect 2413 843 2417 844
rect 2367 838 2391 842
rect 2397 839 2410 843
rect 2367 834 2371 838
rect 2366 833 2371 834
rect 2401 837 2410 839
rect 2401 835 2403 837
rect 2370 829 2371 833
rect 2375 829 2376 833
rect 2380 829 2392 833
rect 2397 830 2403 835
rect 2366 828 2371 829
rect 2367 825 2371 828
rect 2367 824 2384 825
rect 2367 821 2379 824
rect 2378 820 2379 821
rect 2383 820 2384 824
rect 2388 822 2392 829
rect 2413 827 2417 839
rect 2442 837 2446 846
rect 2482 847 2483 851
rect 2487 847 2488 851
rect 2545 847 2546 851
rect 2550 847 2564 851
rect 2471 842 2475 844
rect 2497 843 2501 844
rect 2444 833 2446 837
rect 2451 838 2475 842
rect 2481 839 2494 843
rect 2451 834 2455 838
rect 2405 824 2417 827
rect 2388 820 2405 822
rect 2409 823 2417 824
rect 2388 818 2409 820
rect 2413 818 2418 819
rect 2358 813 2369 817
rect 2373 813 2374 817
rect 2388 814 2392 818
rect 2381 810 2392 814
rect 2417 814 2418 818
rect 2413 811 2418 814
rect 2442 817 2446 833
rect 2450 833 2455 834
rect 2485 837 2494 839
rect 2485 835 2487 837
rect 2454 829 2455 833
rect 2459 829 2460 833
rect 2464 829 2476 833
rect 2481 830 2487 835
rect 2450 828 2455 829
rect 2451 825 2455 828
rect 2451 824 2468 825
rect 2451 821 2463 824
rect 2462 820 2463 821
rect 2467 820 2468 824
rect 2472 822 2476 829
rect 2497 827 2501 839
rect 2544 842 2557 843
rect 2544 838 2549 842
rect 2553 838 2557 842
rect 2544 836 2548 838
rect 2489 824 2501 827
rect 2472 820 2489 822
rect 2493 823 2501 824
rect 2560 834 2564 847
rect 2568 848 2580 851
rect 2568 845 2575 848
rect 2579 844 2580 848
rect 2575 843 2580 844
rect 2576 838 2580 843
rect 2472 818 2493 820
rect 2497 818 2502 819
rect 2507 818 2510 832
rect 2544 829 2548 832
rect 2554 830 2568 834
rect 2572 830 2573 834
rect 2554 825 2560 830
rect 2576 826 2580 834
rect 2575 825 2580 826
rect 2442 813 2453 817
rect 2457 813 2458 817
rect 2472 814 2476 818
rect 2395 810 2399 811
rect 2381 809 2385 810
rect 2358 805 2359 809
rect 2363 805 2385 809
rect 2395 803 2399 806
rect 2406 810 2418 811
rect 2406 806 2409 810
rect 2413 806 2418 810
rect 2465 810 2476 814
rect 2501 815 2510 818
rect 2545 821 2549 822
rect 2554 821 2555 825
rect 2559 821 2560 825
rect 2564 821 2565 825
rect 2569 821 2572 825
rect 2501 814 2502 815
rect 2497 811 2502 814
rect 2479 810 2483 811
rect 2465 809 2469 810
rect 2406 805 2418 806
rect 2442 805 2443 809
rect 2447 805 2469 809
rect 2308 796 2314 800
rect 2318 796 2328 800
rect 2332 796 2342 800
rect 2346 796 2379 800
rect 2383 799 2395 800
rect 2479 803 2483 806
rect 2490 805 2502 811
rect 2399 799 2463 800
rect 2383 796 2463 799
rect 2467 799 2479 800
rect 2545 800 2549 817
rect 2559 811 2565 818
rect 2552 810 2565 811
rect 2556 806 2558 810
rect 2562 806 2565 810
rect 2552 805 2565 806
rect 2568 800 2572 821
rect 2579 821 2580 825
rect 2575 820 2580 821
rect 2576 813 2580 820
rect 2610 800 2614 911
rect 2678 910 2683 913
rect 2678 906 2679 910
rect 2678 905 2683 906
rect 2692 910 2698 914
rect 2702 910 2706 911
rect 2714 910 2737 914
rect 2741 910 2754 914
rect 2678 883 2682 905
rect 2692 901 2696 910
rect 2692 896 2696 897
rect 2699 902 2706 906
rect 2709 902 2747 906
rect 2699 891 2703 902
rect 2709 899 2714 902
rect 2706 898 2714 899
rect 2742 898 2746 902
rect 2710 894 2714 898
rect 2722 894 2725 898
rect 2729 894 2732 898
rect 2736 894 2739 898
rect 2706 893 2714 894
rect 2685 887 2686 891
rect 2690 889 2703 891
rect 2719 889 2723 890
rect 2690 887 2709 889
rect 2699 885 2709 887
rect 2713 885 2714 889
rect 2726 885 2730 894
rect 2742 893 2746 894
rect 2750 899 2754 910
rect 2761 910 2763 914
rect 2757 907 2763 910
rect 2761 903 2763 907
rect 2757 902 2763 903
rect 2750 898 2756 899
rect 2750 894 2752 898
rect 2750 893 2756 894
rect 2750 890 2754 893
rect 2734 886 2754 890
rect 2678 882 2683 883
rect 2678 878 2679 882
rect 2719 882 2723 885
rect 2734 882 2738 886
rect 2759 882 2763 902
rect 2678 877 2683 878
rect 2689 878 2693 879
rect 2698 877 2699 881
rect 2703 878 2719 881
rect 2728 878 2729 882
rect 2733 878 2738 882
rect 2741 878 2757 882
rect 2761 878 2763 882
rect 2703 877 2723 878
rect 2689 872 2693 874
rect 2745 872 2746 875
rect 2674 871 2746 872
rect 2750 872 2751 875
rect 2788 874 2791 918
rect 2811 916 2812 920
rect 2816 918 2824 920
rect 2827 918 2842 922
rect 2846 918 2847 922
rect 2811 915 2816 916
rect 2811 885 2815 915
rect 2827 914 2831 918
rect 2819 910 2831 914
rect 2835 912 2852 915
rect 2819 899 2823 910
rect 2835 906 2839 912
rect 2826 902 2829 906
rect 2833 902 2839 906
rect 2819 891 2823 895
rect 2834 894 2839 898
rect 2843 893 2847 903
rect 2878 898 2881 924
rect 2970 913 2975 933
rect 2819 887 2836 891
rect 2872 887 2951 890
rect 2811 884 2816 885
rect 2832 884 2836 887
rect 2811 880 2812 884
rect 2811 877 2816 880
rect 2821 880 2822 884
rect 2826 880 2827 884
rect 2750 871 2774 872
rect 2674 866 2774 871
rect 2821 872 2827 880
rect 2832 879 2836 880
rect 2841 880 2842 884
rect 2846 880 2847 884
rect 2841 872 2847 880
rect 2854 878 2951 881
rect 2955 878 2957 881
rect 2807 868 2813 872
rect 2817 868 2841 872
rect 2845 868 2851 872
rect 2807 866 2851 868
rect 2668 864 2941 866
rect 2483 799 2546 800
rect 2467 796 2546 799
rect 2550 796 2560 800
rect 2564 796 2574 800
rect 2578 796 2614 800
rect 2308 792 2614 796
rect 2308 786 2309 792
rect 2315 786 2614 792
rect 2308 784 2614 786
rect 2307 782 2614 784
rect 2634 862 2941 864
rect 2634 859 2692 862
rect 2307 780 2613 782
rect 2307 776 2343 780
rect 2347 776 2357 780
rect 2361 776 2371 780
rect 2375 777 2454 780
rect 2375 776 2438 777
rect 2233 733 2247 737
rect 2251 733 2252 737
rect 2279 736 2280 741
rect 1984 724 1987 728
rect 1991 724 1997 728
rect 2001 724 2065 728
rect 2069 724 2118 728
rect 2122 724 2149 728
rect 2153 724 2202 728
rect 2206 724 2219 728
rect 2223 724 2229 728
rect 2233 724 2257 728
rect 1984 723 2257 724
rect 1970 720 2257 723
rect 1970 716 2070 720
rect 1970 715 1994 716
rect 1993 712 1994 715
rect 1998 715 2070 716
rect 2074 718 2118 720
rect 1998 712 1999 715
rect 2051 713 2055 715
rect 2074 714 2080 718
rect 2084 714 2108 718
rect 2112 714 2118 718
rect 2021 709 2041 710
rect 1950 653 1955 673
rect 1981 705 1983 709
rect 1987 705 1994 709
rect 1998 705 2003 709
rect 2006 705 2011 709
rect 2015 705 2016 709
rect 2025 706 2041 709
rect 2045 706 2046 710
rect 2051 708 2055 709
rect 2061 709 2066 710
rect 1981 685 1985 705
rect 2006 701 2010 705
rect 2021 702 2025 705
rect 2065 705 2066 709
rect 2061 704 2066 705
rect 1990 697 2010 701
rect 1990 694 1994 697
rect 1988 693 1994 694
rect 1992 689 1994 693
rect 1988 688 1994 689
rect 1981 684 1987 685
rect 1981 680 1983 684
rect 1981 677 1987 680
rect 1981 673 1983 677
rect 1990 677 1994 688
rect 1998 693 2002 694
rect 2014 693 2018 702
rect 2030 698 2031 702
rect 2035 700 2045 702
rect 2035 698 2054 700
rect 2021 697 2025 698
rect 2041 696 2054 698
rect 2058 696 2059 700
rect 2030 693 2038 694
rect 2005 689 2008 693
rect 2012 689 2015 693
rect 2019 689 2020 693
rect 2030 689 2034 693
rect 1998 685 2002 689
rect 2030 688 2038 689
rect 2030 685 2035 688
rect 2041 685 2045 696
rect 1997 681 2035 685
rect 2038 681 2045 685
rect 2048 690 2052 691
rect 2048 677 2052 686
rect 2062 682 2066 704
rect 2078 706 2084 714
rect 2078 702 2079 706
rect 2083 702 2084 706
rect 2089 706 2093 707
rect 2098 706 2104 714
rect 2098 702 2099 706
rect 2103 702 2104 706
rect 2109 706 2114 709
rect 2113 702 2114 706
rect 2089 699 2093 702
rect 2109 701 2114 702
rect 2089 695 2106 699
rect 1990 673 2003 677
rect 2007 673 2030 677
rect 2038 676 2042 677
rect 2046 673 2052 677
rect 2061 681 2066 682
rect 2065 677 2066 681
rect 2078 683 2082 693
rect 2086 688 2091 692
rect 2102 691 2106 695
rect 2086 680 2092 684
rect 2096 680 2099 684
rect 2061 674 2066 677
rect 1981 672 1987 673
rect 2003 670 2007 673
rect 1992 665 1993 669
rect 1997 665 1998 669
rect 2026 669 2050 673
rect 2065 670 2066 674
rect 2086 674 2090 680
rect 2102 676 2106 687
rect 2073 671 2090 674
rect 2094 672 2106 676
rect 2110 696 2114 701
rect 2110 690 2229 696
rect 2061 669 2066 670
rect 2003 665 2007 666
rect 2014 665 2015 669
rect 2019 665 2020 669
rect 2053 668 2066 669
rect 2094 668 2098 672
rect 2110 671 2114 690
rect 2226 684 2229 690
rect 2109 670 2114 671
rect 2053 667 2067 668
rect 2053 665 2065 667
rect 1992 662 1998 665
rect 1992 659 1993 662
rect 1970 658 1993 659
rect 1997 659 1998 662
rect 2014 662 2020 665
rect 2064 663 2065 665
rect 2069 663 2071 666
rect 2078 664 2079 668
rect 2083 664 2098 668
rect 2101 666 2109 668
rect 2113 666 2114 670
rect 2101 664 2114 666
rect 2251 667 2256 720
rect 2295 718 2300 761
rect 2251 662 2293 667
rect 2298 662 2299 667
rect 2307 665 2311 776
rect 2341 756 2345 763
rect 2341 755 2346 756
rect 2341 751 2342 755
rect 2349 755 2353 776
rect 2356 770 2369 771
rect 2356 766 2359 770
rect 2363 766 2365 770
rect 2356 765 2369 766
rect 2356 758 2362 765
rect 2372 759 2376 776
rect 2442 776 2454 777
rect 2458 777 2538 780
rect 2458 776 2522 777
rect 2419 765 2431 771
rect 2438 770 2442 773
rect 2526 776 2538 777
rect 2542 776 2575 780
rect 2579 776 2589 780
rect 2593 776 2603 780
rect 2607 776 2613 780
rect 2452 767 2474 771
rect 2478 767 2479 771
rect 2452 766 2456 767
rect 2438 765 2442 766
rect 2419 762 2424 765
rect 2419 761 2420 762
rect 2411 758 2420 761
rect 2445 762 2456 766
rect 2445 758 2449 762
rect 2463 759 2464 763
rect 2468 759 2479 763
rect 2349 751 2352 755
rect 2356 751 2357 755
rect 2361 751 2362 755
rect 2366 751 2367 755
rect 2372 754 2376 755
rect 2341 750 2346 751
rect 2341 742 2345 750
rect 2361 746 2367 751
rect 2348 742 2349 746
rect 2353 742 2367 746
rect 2373 744 2377 747
rect 2341 733 2345 738
rect 2341 732 2346 733
rect 2341 728 2342 732
rect 2346 728 2353 731
rect 2341 725 2353 728
rect 2357 729 2361 742
rect 2373 738 2377 740
rect 2364 734 2368 738
rect 2372 734 2377 738
rect 2364 733 2377 734
rect 2401 736 2405 750
rect 2411 744 2414 758
rect 2419 757 2424 758
rect 2428 756 2449 758
rect 2420 752 2428 753
rect 2432 754 2449 756
rect 2420 749 2432 752
rect 2420 737 2424 749
rect 2445 747 2449 754
rect 2453 752 2454 756
rect 2458 755 2459 756
rect 2458 752 2470 755
rect 2453 751 2470 752
rect 2466 748 2470 751
rect 2466 747 2471 748
rect 2434 741 2440 746
rect 2445 743 2457 747
rect 2461 743 2462 747
rect 2466 743 2467 747
rect 2434 739 2436 741
rect 2427 737 2436 739
rect 2466 742 2471 743
rect 2475 743 2479 759
rect 2466 738 2470 742
rect 2427 733 2440 737
rect 2446 734 2470 738
rect 2475 739 2477 743
rect 2420 732 2424 733
rect 2446 732 2450 734
rect 2357 725 2371 729
rect 2375 725 2376 729
rect 2433 725 2434 729
rect 2438 725 2439 729
rect 2475 730 2479 739
rect 2446 727 2450 728
rect 2455 726 2456 730
rect 2460 726 2479 730
rect 2489 728 2492 767
rect 2503 770 2515 771
rect 2503 766 2508 770
rect 2512 766 2515 770
rect 2503 765 2515 766
rect 2522 770 2526 773
rect 2536 767 2558 771
rect 2562 767 2563 771
rect 2536 766 2540 767
rect 2522 765 2526 766
rect 2503 762 2508 765
rect 2503 758 2504 762
rect 2529 762 2540 766
rect 2529 758 2533 762
rect 2547 759 2548 763
rect 2552 759 2563 763
rect 2503 757 2508 758
rect 2512 756 2533 758
rect 2504 752 2512 753
rect 2516 754 2533 756
rect 2504 749 2516 752
rect 2504 737 2508 749
rect 2529 747 2533 754
rect 2537 752 2538 756
rect 2542 755 2543 756
rect 2542 752 2554 755
rect 2537 751 2554 752
rect 2550 748 2554 751
rect 2559 752 2563 759
rect 2573 756 2577 763
rect 2573 755 2578 756
rect 2559 749 2566 752
rect 2573 751 2574 755
rect 2581 755 2585 776
rect 2588 770 2601 771
rect 2588 766 2591 770
rect 2595 766 2597 770
rect 2588 765 2601 766
rect 2588 758 2594 765
rect 2604 759 2608 776
rect 2581 751 2584 755
rect 2588 751 2589 755
rect 2593 751 2594 755
rect 2598 751 2599 755
rect 2604 754 2608 755
rect 2573 750 2578 751
rect 2550 747 2555 748
rect 2518 741 2524 746
rect 2529 743 2541 747
rect 2545 743 2546 747
rect 2550 743 2551 747
rect 2518 739 2520 741
rect 2511 737 2520 739
rect 2550 742 2555 743
rect 2550 738 2554 742
rect 2511 733 2524 737
rect 2530 734 2554 738
rect 2504 732 2508 733
rect 2530 732 2534 734
rect 2433 720 2439 725
rect 2517 725 2518 729
rect 2522 725 2523 729
rect 2559 730 2563 749
rect 2573 742 2577 750
rect 2593 746 2599 751
rect 2580 742 2581 746
rect 2585 742 2599 746
rect 2605 745 2609 747
rect 2530 727 2534 728
rect 2539 726 2540 730
rect 2544 726 2563 730
rect 2567 739 2577 742
rect 2567 727 2570 739
rect 2489 723 2492 724
rect 2517 720 2523 725
rect 2573 733 2577 739
rect 2573 732 2578 733
rect 2573 728 2574 732
rect 2578 728 2585 731
rect 2573 725 2585 728
rect 2589 729 2593 742
rect 2634 743 2640 859
rect 2668 858 2692 859
rect 2696 858 2702 862
rect 2706 858 2719 862
rect 2723 858 2772 862
rect 2776 858 2803 862
rect 2807 858 2856 862
rect 2860 858 2924 862
rect 2928 858 2934 862
rect 2938 858 2941 862
rect 2673 849 2674 853
rect 2678 849 2692 853
rect 2672 844 2685 845
rect 2672 840 2677 844
rect 2681 840 2685 844
rect 2672 837 2676 840
rect 2688 836 2692 849
rect 2696 850 2708 853
rect 2696 847 2703 850
rect 2707 846 2708 850
rect 2703 845 2708 846
rect 2704 839 2708 845
rect 2758 853 2764 858
rect 2711 839 2714 851
rect 2704 836 2714 839
rect 2718 848 2737 852
rect 2741 848 2742 852
rect 2747 850 2751 851
rect 2672 831 2676 833
rect 2682 832 2696 836
rect 2700 832 2701 836
rect 2682 827 2688 832
rect 2704 828 2708 836
rect 2703 827 2708 828
rect 2718 827 2722 848
rect 2758 849 2759 853
rect 2763 849 2764 853
rect 2786 851 2791 855
rect 2842 853 2848 858
rect 2747 844 2751 846
rect 2773 845 2777 846
rect 2727 840 2751 844
rect 2757 841 2770 845
rect 2727 836 2731 840
rect 2726 835 2731 836
rect 2761 839 2770 841
rect 2761 837 2763 839
rect 2730 831 2731 835
rect 2735 831 2736 835
rect 2740 831 2752 835
rect 2757 832 2763 837
rect 2726 830 2731 831
rect 2673 823 2677 824
rect 2682 823 2683 827
rect 2687 823 2688 827
rect 2692 823 2693 827
rect 2697 823 2700 827
rect 2673 802 2677 819
rect 2687 813 2693 820
rect 2680 812 2693 813
rect 2684 808 2686 812
rect 2690 808 2693 812
rect 2680 807 2693 808
rect 2696 802 2700 823
rect 2707 823 2708 827
rect 2716 823 2722 827
rect 2727 827 2731 830
rect 2727 826 2744 827
rect 2727 823 2739 826
rect 2703 822 2708 823
rect 2704 815 2708 822
rect 2718 819 2722 823
rect 2738 822 2739 823
rect 2743 822 2744 826
rect 2748 824 2752 831
rect 2773 829 2777 841
rect 2765 826 2777 829
rect 2788 828 2791 851
rect 2802 848 2821 852
rect 2825 848 2826 852
rect 2831 850 2835 851
rect 2802 839 2806 848
rect 2842 849 2843 853
rect 2847 849 2848 853
rect 2905 849 2906 853
rect 2910 849 2924 853
rect 2831 844 2835 846
rect 2857 845 2861 846
rect 2804 835 2806 839
rect 2811 840 2835 844
rect 2841 841 2854 845
rect 2811 836 2815 840
rect 2748 822 2765 824
rect 2769 825 2777 826
rect 2748 820 2769 822
rect 2773 820 2778 821
rect 2718 815 2729 819
rect 2733 815 2734 819
rect 2748 816 2752 820
rect 2741 812 2752 816
rect 2777 816 2778 820
rect 2773 813 2778 816
rect 2802 819 2806 835
rect 2810 835 2815 836
rect 2845 839 2854 841
rect 2845 837 2847 839
rect 2814 831 2815 835
rect 2819 831 2820 835
rect 2824 831 2836 835
rect 2841 832 2847 837
rect 2810 830 2815 831
rect 2811 827 2815 830
rect 2811 826 2828 827
rect 2811 823 2823 826
rect 2822 822 2823 823
rect 2827 822 2828 826
rect 2832 824 2836 831
rect 2857 829 2861 841
rect 2904 844 2917 845
rect 2904 840 2909 844
rect 2913 840 2917 844
rect 2904 838 2908 840
rect 2849 826 2861 829
rect 2832 822 2849 824
rect 2853 825 2861 826
rect 2920 836 2924 849
rect 2928 850 2940 853
rect 2928 847 2935 850
rect 2939 846 2940 850
rect 2935 845 2940 846
rect 2936 840 2940 845
rect 2832 820 2853 822
rect 2857 820 2862 821
rect 2867 820 2870 834
rect 2904 831 2908 834
rect 2914 832 2928 836
rect 2932 832 2933 836
rect 2914 827 2920 832
rect 2936 828 2940 836
rect 2935 827 2940 828
rect 2802 815 2813 819
rect 2817 815 2818 819
rect 2832 816 2836 820
rect 2755 812 2759 813
rect 2741 811 2745 812
rect 2718 807 2719 811
rect 2723 807 2745 811
rect 2755 805 2759 808
rect 2766 812 2778 813
rect 2766 808 2769 812
rect 2773 808 2778 812
rect 2825 812 2836 816
rect 2861 817 2870 820
rect 2905 823 2909 824
rect 2914 823 2915 827
rect 2919 823 2920 827
rect 2924 823 2925 827
rect 2929 823 2932 827
rect 2861 816 2862 817
rect 2857 813 2862 816
rect 2839 812 2843 813
rect 2825 811 2829 812
rect 2766 807 2778 808
rect 2802 807 2803 811
rect 2807 807 2829 811
rect 2668 798 2674 802
rect 2678 798 2688 802
rect 2692 798 2702 802
rect 2706 798 2739 802
rect 2743 801 2755 802
rect 2839 805 2843 808
rect 2850 807 2862 813
rect 2759 801 2823 802
rect 2743 798 2823 801
rect 2827 801 2839 802
rect 2905 802 2909 819
rect 2919 813 2925 820
rect 2912 812 2925 813
rect 2916 808 2918 812
rect 2922 808 2925 812
rect 2912 807 2925 808
rect 2928 802 2932 823
rect 2939 823 2940 827
rect 2935 822 2940 823
rect 2936 815 2940 822
rect 2970 802 2974 913
rect 2843 801 2906 802
rect 2827 798 2906 801
rect 2910 798 2920 802
rect 2924 798 2934 802
rect 2938 798 2974 802
rect 2668 786 2974 798
rect 2605 738 2609 741
rect 2596 734 2600 738
rect 2604 734 2609 738
rect 2596 733 2609 734
rect 2632 736 2633 741
rect 2639 738 2640 743
rect 2667 784 2974 786
rect 2667 782 2973 784
rect 2667 778 2703 782
rect 2707 778 2717 782
rect 2721 778 2731 782
rect 2735 779 2814 782
rect 2735 778 2798 779
rect 2589 725 2603 729
rect 2607 725 2608 729
rect 2340 716 2343 720
rect 2347 716 2353 720
rect 2357 716 2421 720
rect 2425 716 2474 720
rect 2478 716 2505 720
rect 2509 716 2558 720
rect 2562 716 2575 720
rect 2579 716 2585 720
rect 2589 718 2613 720
rect 2632 718 2638 736
rect 2589 716 2643 718
rect 2323 714 2643 716
rect 2326 713 2643 714
rect 2326 712 2613 713
rect 2326 706 2404 712
rect 2430 710 2474 712
rect 2430 706 2436 710
rect 2440 706 2464 710
rect 2468 706 2474 710
rect 2343 666 2348 706
rect 2434 698 2440 706
rect 2434 694 2435 698
rect 2439 694 2440 698
rect 2445 698 2449 699
rect 2454 698 2460 706
rect 2454 694 2455 698
rect 2459 694 2460 698
rect 2465 698 2470 701
rect 2469 694 2470 698
rect 2445 691 2449 694
rect 2465 693 2470 694
rect 2445 687 2462 691
rect 2014 659 2015 662
rect 1997 658 2015 659
rect 2019 659 2020 662
rect 2049 659 2050 662
rect 2019 658 2050 659
rect 2054 659 2055 662
rect 2054 658 2070 659
rect 2096 658 2097 661
rect 1970 656 2070 658
rect 1968 653 2070 656
rect 2074 657 2097 658
rect 2101 658 2102 661
rect 2101 657 2108 658
rect 2074 654 2108 657
rect 2112 654 2118 658
rect 2074 653 2118 654
rect 1950 650 2118 653
rect 1950 649 2074 650
rect 1922 640 1953 644
rect 1922 637 1954 640
rect 1902 522 1905 633
rect 1914 611 1919 612
rect 1914 564 1919 606
rect 1929 574 1934 619
rect 1914 553 1920 564
rect 1885 478 1892 493
rect 1885 329 1891 478
rect 1915 428 1920 553
rect 1945 546 1954 637
rect 1952 541 1954 546
rect 1982 481 1987 649
rect 2268 645 2272 662
rect 2306 645 2311 665
rect 2402 664 2405 685
rect 2434 675 2438 685
rect 2442 680 2447 684
rect 2458 683 2462 687
rect 2442 672 2448 676
rect 2452 672 2455 676
rect 2442 666 2446 672
rect 2458 668 2462 679
rect 2429 663 2446 666
rect 2450 664 2462 668
rect 2466 689 2470 693
rect 2489 689 2492 702
rect 2466 686 2492 689
rect 2450 660 2454 664
rect 2466 663 2470 686
rect 2667 667 2671 778
rect 2701 758 2705 765
rect 2701 757 2706 758
rect 2701 753 2702 757
rect 2709 757 2713 778
rect 2716 772 2729 773
rect 2716 768 2719 772
rect 2723 768 2725 772
rect 2716 767 2729 768
rect 2716 760 2722 767
rect 2732 761 2736 778
rect 2802 778 2814 779
rect 2818 779 2898 782
rect 2818 778 2882 779
rect 2779 767 2791 773
rect 2798 772 2802 775
rect 2886 778 2898 779
rect 2902 778 2935 782
rect 2939 778 2949 782
rect 2953 778 2963 782
rect 2967 778 2973 782
rect 2812 769 2834 773
rect 2838 769 2839 773
rect 2812 768 2816 769
rect 2798 767 2802 768
rect 2779 764 2784 767
rect 2779 763 2780 764
rect 2709 753 2712 757
rect 2716 753 2717 757
rect 2721 753 2722 757
rect 2726 753 2727 757
rect 2732 756 2736 757
rect 2771 760 2780 763
rect 2805 764 2816 768
rect 2805 760 2809 764
rect 2823 761 2824 765
rect 2828 761 2839 765
rect 2701 752 2706 753
rect 2701 744 2705 752
rect 2721 748 2727 753
rect 2708 744 2709 748
rect 2713 744 2727 748
rect 2733 746 2737 749
rect 2701 735 2705 740
rect 2701 734 2706 735
rect 2701 730 2702 734
rect 2706 730 2713 733
rect 2701 727 2713 730
rect 2717 731 2721 744
rect 2733 740 2737 742
rect 2724 736 2728 740
rect 2732 736 2737 740
rect 2724 735 2737 736
rect 2752 735 2755 752
rect 2771 746 2774 760
rect 2779 759 2784 760
rect 2788 758 2809 760
rect 2780 754 2788 755
rect 2792 756 2809 758
rect 2780 751 2792 754
rect 2780 739 2784 751
rect 2805 749 2809 756
rect 2813 754 2814 758
rect 2818 757 2819 758
rect 2818 754 2830 757
rect 2813 753 2830 754
rect 2826 750 2830 753
rect 2826 749 2831 750
rect 2794 743 2800 748
rect 2805 745 2817 749
rect 2821 745 2822 749
rect 2826 745 2827 749
rect 2794 741 2796 743
rect 2787 739 2796 741
rect 2826 744 2831 745
rect 2835 745 2839 761
rect 2826 740 2830 744
rect 2787 735 2800 739
rect 2806 736 2830 740
rect 2835 741 2837 745
rect 2780 734 2784 735
rect 2806 734 2810 736
rect 2717 727 2731 731
rect 2735 727 2736 731
rect 2793 727 2794 731
rect 2798 727 2799 731
rect 2835 732 2839 741
rect 2806 729 2810 730
rect 2815 728 2816 732
rect 2820 728 2839 732
rect 2849 730 2852 769
rect 2863 772 2875 773
rect 2863 768 2868 772
rect 2872 768 2875 772
rect 2863 767 2875 768
rect 2882 772 2886 775
rect 2896 769 2918 773
rect 2922 769 2923 773
rect 2896 768 2900 769
rect 2882 767 2886 768
rect 2863 764 2868 767
rect 2863 760 2864 764
rect 2889 764 2900 768
rect 2889 760 2893 764
rect 2907 761 2908 765
rect 2912 761 2923 765
rect 2863 759 2868 760
rect 2872 758 2893 760
rect 2864 754 2872 755
rect 2876 756 2893 758
rect 2864 751 2876 754
rect 2864 739 2868 751
rect 2889 749 2893 756
rect 2897 754 2898 758
rect 2902 757 2903 758
rect 2902 754 2914 757
rect 2897 753 2914 754
rect 2910 750 2914 753
rect 2919 754 2923 761
rect 2933 758 2937 765
rect 2933 757 2938 758
rect 2910 749 2915 750
rect 2878 743 2884 748
rect 2889 745 2901 749
rect 2905 745 2906 749
rect 2910 745 2911 749
rect 2878 741 2880 743
rect 2871 739 2880 741
rect 2910 744 2915 745
rect 2919 749 2925 754
rect 2933 753 2934 757
rect 2941 757 2945 778
rect 2948 772 2961 773
rect 2948 768 2951 772
rect 2955 768 2957 772
rect 2948 767 2961 768
rect 2948 760 2954 767
rect 2964 761 2968 778
rect 2941 753 2944 757
rect 2948 753 2949 757
rect 2953 753 2954 757
rect 2958 753 2959 757
rect 2964 756 2968 757
rect 2933 752 2938 753
rect 2910 740 2914 744
rect 2871 735 2884 739
rect 2890 736 2914 740
rect 2864 734 2868 735
rect 2890 734 2894 736
rect 2793 722 2799 727
rect 2877 727 2878 731
rect 2882 727 2883 731
rect 2919 732 2923 749
rect 2933 744 2937 752
rect 2953 748 2959 753
rect 2940 744 2941 748
rect 2945 744 2959 748
rect 2890 729 2894 730
rect 2899 728 2900 732
rect 2904 728 2923 732
rect 2927 741 2937 744
rect 2927 729 2930 741
rect 2849 725 2852 726
rect 2877 722 2883 727
rect 2933 735 2937 741
rect 2933 734 2938 735
rect 2933 730 2934 734
rect 2938 730 2945 733
rect 2933 727 2945 730
rect 2949 731 2953 744
rect 2965 740 2969 743
rect 2956 736 2960 740
rect 2964 736 2969 740
rect 2956 735 2969 736
rect 2949 727 2963 731
rect 2967 727 2968 731
rect 2700 718 2703 722
rect 2707 718 2713 722
rect 2717 718 2781 722
rect 2785 718 2834 722
rect 2838 718 2865 722
rect 2869 718 2918 722
rect 2922 718 2935 722
rect 2939 718 2945 722
rect 2949 718 2973 722
rect 2683 716 2973 718
rect 2686 714 2973 716
rect 2686 708 2764 714
rect 2790 712 2834 714
rect 2790 708 2796 712
rect 2800 708 2824 712
rect 2828 708 2834 712
rect 2794 700 2800 708
rect 2794 696 2795 700
rect 2799 696 2800 700
rect 2805 700 2809 701
rect 2814 700 2820 708
rect 2814 696 2815 700
rect 2819 696 2820 700
rect 2825 700 2830 703
rect 2829 696 2830 700
rect 2465 662 2470 663
rect 2434 656 2435 660
rect 2439 656 2454 660
rect 2457 658 2465 660
rect 2469 658 2470 662
rect 2457 656 2470 658
rect 2452 650 2453 653
rect 2430 649 2453 650
rect 2457 650 2458 653
rect 2457 649 2464 650
rect 2430 646 2464 649
rect 2468 648 2474 650
rect 2666 648 2671 667
rect 2754 668 2757 694
rect 2805 693 2809 696
rect 2825 695 2830 696
rect 2805 689 2822 693
rect 2763 667 2766 680
rect 2794 677 2798 687
rect 2802 682 2807 686
rect 2818 685 2822 689
rect 2802 674 2808 678
rect 2812 674 2815 678
rect 2802 668 2806 674
rect 2818 670 2822 681
rect 2789 665 2806 668
rect 2810 666 2822 670
rect 2826 691 2830 695
rect 2849 691 2852 704
rect 2826 688 2852 691
rect 2810 662 2814 666
rect 2826 665 2830 688
rect 2825 664 2830 665
rect 2794 658 2795 662
rect 2799 658 2814 662
rect 2817 660 2825 662
rect 2829 660 2830 664
rect 2817 658 2830 660
rect 2812 652 2813 655
rect 2468 647 2671 648
rect 2790 651 2813 652
rect 2817 652 2818 655
rect 2817 651 2824 652
rect 2790 648 2824 651
rect 2828 648 2834 652
rect 2790 647 2834 648
rect 2468 646 2834 647
rect 2430 645 2834 646
rect 2306 644 2834 645
rect 2306 643 2790 644
rect 2306 642 2670 643
rect 2306 641 2430 642
rect 2013 636 2019 639
rect 2033 629 2036 633
rect 1998 628 2037 629
rect 1994 626 2037 628
rect 2064 590 2067 634
rect 2623 625 2957 628
rect 2064 587 2959 590
rect 2035 504 2038 585
rect 2262 571 2267 573
rect 2266 567 2267 571
rect 2034 500 2251 504
rect 2247 495 2251 500
rect 2262 482 2267 567
rect 1986 476 1987 481
rect 2202 477 2267 482
rect 1952 465 2393 469
rect 1952 443 1956 465
rect 1980 458 1981 462
rect 1902 414 1962 418
rect 1980 377 1984 458
rect 2034 456 2035 459
rect 2034 455 2197 456
rect 2029 454 2197 455
rect 2250 456 2443 457
rect 2449 456 2493 458
rect 2202 455 2493 456
rect 2542 455 2586 458
rect 2629 457 2673 458
rect 2629 455 2681 457
rect 2202 454 2681 455
rect 2029 452 2455 454
rect 2029 448 2053 452
rect 2057 448 2063 452
rect 2067 448 2140 452
rect 2144 448 2150 452
rect 2154 448 2233 452
rect 2237 448 2243 452
rect 2247 451 2455 452
rect 2247 448 2253 451
rect 2449 450 2455 451
rect 2459 450 2465 454
rect 2469 451 2548 454
rect 2469 450 2493 451
rect 2542 450 2548 451
rect 2552 450 2558 454
rect 2562 451 2635 454
rect 2562 450 2586 451
rect 2629 450 2635 451
rect 2639 450 2645 454
rect 2649 451 2681 454
rect 2649 450 2673 451
rect 2033 438 2034 442
rect 2038 438 2053 442
rect 1999 432 2029 435
rect 2033 431 2045 435
rect 2040 426 2045 431
rect 2049 434 2053 438
rect 2057 440 2069 443
rect 2057 437 2064 440
rect 2068 436 2069 440
rect 2120 438 2121 442
rect 2125 438 2140 442
rect 2064 435 2069 436
rect 2049 430 2061 434
rect 2057 426 2061 430
rect 2040 422 2047 426
rect 2051 422 2054 426
rect 2033 409 2037 418
rect 2041 414 2046 418
rect 2057 411 2061 422
rect 2065 421 2069 435
rect 2121 431 2132 435
rect 2127 426 2132 431
rect 2136 434 2140 438
rect 2144 440 2156 443
rect 2144 437 2151 440
rect 2155 436 2156 440
rect 2213 438 2214 442
rect 2218 438 2233 442
rect 2151 435 2156 436
rect 2136 430 2148 434
rect 2144 426 2148 430
rect 2127 422 2134 426
rect 2138 422 2141 426
rect 2065 418 2094 421
rect 2065 417 2069 418
rect 2026 405 2037 409
rect 2044 409 2061 411
rect 2048 407 2061 409
rect 2064 416 2069 417
rect 2068 412 2069 416
rect 2064 409 2069 412
rect 2044 402 2048 405
rect 2068 405 2069 409
rect 2064 404 2069 405
rect 2033 398 2034 402
rect 2038 398 2039 402
rect 2033 392 2039 398
rect 2044 397 2048 398
rect 2053 400 2054 404
rect 2058 400 2059 404
rect 2053 392 2059 400
rect 2029 388 2063 392
rect 2067 388 2073 392
rect 2029 384 2073 388
rect 2030 377 2034 384
rect 2090 382 2094 418
rect 2120 408 2124 418
rect 2128 414 2133 418
rect 2144 411 2148 422
rect 2152 417 2156 435
rect 2214 431 2225 435
rect 2220 426 2225 431
rect 2229 434 2233 438
rect 2237 440 2249 443
rect 2453 442 2465 445
rect 2237 437 2244 440
rect 2248 436 2249 440
rect 2262 436 2434 440
rect 2439 436 2440 440
rect 2453 438 2454 442
rect 2458 439 2465 442
rect 2469 440 2484 444
rect 2488 440 2489 444
rect 2546 442 2558 445
rect 2453 437 2458 438
rect 2244 435 2249 436
rect 2229 430 2241 434
rect 2237 426 2241 430
rect 2220 422 2227 426
rect 2231 422 2234 426
rect 2117 405 2124 408
rect 2131 409 2148 411
rect 2135 407 2148 409
rect 2151 416 2156 417
rect 2155 412 2156 416
rect 2151 409 2156 412
rect 2131 402 2135 405
rect 2155 407 2156 409
rect 2155 405 2162 407
rect 2151 404 2162 405
rect 2213 408 2217 418
rect 2221 414 2226 418
rect 2237 411 2241 422
rect 2245 431 2249 435
rect 2245 427 2293 431
rect 2453 430 2457 437
rect 2469 436 2473 440
rect 2546 438 2547 442
rect 2551 439 2558 442
rect 2562 440 2577 444
rect 2581 440 2582 444
rect 2633 442 2645 445
rect 2546 437 2551 438
rect 2245 417 2249 427
rect 2397 426 2457 430
rect 2453 419 2457 426
rect 2461 432 2473 436
rect 2477 434 2488 437
rect 2461 428 2465 432
rect 2477 428 2482 434
rect 2468 424 2471 428
rect 2475 424 2482 428
rect 2546 426 2550 437
rect 2562 436 2566 440
rect 2633 438 2634 442
rect 2638 439 2645 442
rect 2649 440 2664 444
rect 2668 440 2669 444
rect 2633 437 2638 438
rect 2453 418 2458 419
rect 2210 405 2217 408
rect 2224 409 2241 411
rect 2228 407 2241 409
rect 2244 416 2249 417
rect 2248 412 2249 416
rect 2262 414 2435 417
rect 2453 414 2454 418
rect 2244 409 2249 412
rect 2120 398 2121 402
rect 2125 398 2126 402
rect 2120 392 2126 398
rect 2131 397 2135 398
rect 2140 400 2141 404
rect 2145 400 2146 404
rect 2224 402 2228 405
rect 2248 405 2249 409
rect 2453 411 2458 414
rect 2453 407 2454 411
rect 2461 413 2465 424
rect 2523 423 2550 426
rect 2476 416 2481 420
rect 2461 411 2478 413
rect 2461 409 2474 411
rect 2453 406 2458 407
rect 2485 410 2489 420
rect 2523 411 2527 423
rect 2485 407 2492 410
rect 2244 404 2249 405
rect 2140 392 2146 400
rect 2213 398 2214 402
rect 2218 398 2219 402
rect 2213 392 2219 398
rect 2224 397 2228 398
rect 2233 400 2234 404
rect 2238 400 2239 404
rect 2463 402 2464 406
rect 2468 402 2469 406
rect 2233 392 2239 400
rect 2262 396 2436 399
rect 2463 394 2469 402
rect 2474 404 2478 407
rect 2546 419 2550 423
rect 2554 432 2566 436
rect 2570 436 2584 437
rect 2570 434 2581 436
rect 2554 428 2558 432
rect 2570 428 2575 434
rect 2561 424 2564 428
rect 2568 424 2575 428
rect 2546 418 2551 419
rect 2546 414 2547 418
rect 2546 411 2551 414
rect 2546 407 2547 411
rect 2554 413 2558 424
rect 2633 423 2637 437
rect 2649 436 2653 440
rect 2569 416 2574 420
rect 2554 411 2571 413
rect 2554 409 2567 411
rect 2546 406 2551 407
rect 2578 410 2582 420
rect 2611 419 2637 423
rect 2641 432 2653 436
rect 2657 436 2671 437
rect 2657 434 2668 436
rect 2641 428 2645 432
rect 2657 428 2662 434
rect 2648 424 2651 428
rect 2655 424 2662 428
rect 2578 407 2585 410
rect 2597 409 2598 413
rect 2474 399 2478 400
rect 2483 400 2484 404
rect 2488 400 2489 404
rect 2483 394 2489 400
rect 2556 402 2557 406
rect 2561 402 2562 406
rect 2556 394 2562 402
rect 2567 404 2571 407
rect 2567 399 2571 400
rect 2576 400 2577 404
rect 2581 400 2582 404
rect 2576 394 2582 400
rect 2116 388 2150 392
rect 2154 388 2160 392
rect 2116 387 2160 388
rect 2209 388 2243 392
rect 2247 388 2253 392
rect 2116 384 2143 387
rect 2209 384 2253 388
rect 2449 390 2455 394
rect 2459 390 2493 394
rect 2542 390 2548 394
rect 2552 390 2586 394
rect 2449 386 2493 390
rect 2118 377 2122 384
rect 2155 380 2188 383
rect 2209 377 2213 384
rect 2485 382 2489 386
rect 2504 385 2534 388
rect 2542 386 2586 390
rect 2597 389 2601 409
rect 2443 381 2547 382
rect 2443 379 2569 381
rect 2578 379 2582 386
rect 2611 388 2615 419
rect 2633 418 2638 419
rect 2633 414 2634 418
rect 2621 389 2625 409
rect 2633 411 2638 414
rect 2633 407 2634 411
rect 2641 413 2645 424
rect 2656 416 2661 420
rect 2641 411 2658 413
rect 2641 409 2654 411
rect 2633 406 2638 407
rect 2665 411 2669 420
rect 2665 407 2673 411
rect 2643 402 2644 406
rect 2648 402 2649 406
rect 2643 394 2649 402
rect 2654 404 2658 407
rect 2654 399 2658 400
rect 2663 400 2664 404
rect 2668 400 2669 404
rect 2909 401 2913 507
rect 2663 394 2669 400
rect 2629 390 2635 394
rect 2639 390 2673 394
rect 2629 386 2673 390
rect 2667 379 2671 386
rect 2681 379 2883 382
rect 2225 378 2883 379
rect 2225 377 2613 378
rect 1921 376 2148 377
rect 2161 376 2613 377
rect 1921 375 2613 376
rect 1921 373 2286 375
rect 1921 369 1957 373
rect 1961 369 1971 373
rect 1975 369 1985 373
rect 1989 370 2068 373
rect 1989 369 2052 370
rect 1784 289 1878 291
rect 1821 287 1878 289
rect 1873 286 1878 287
rect 1773 271 1784 276
rect 1722 251 1735 253
rect 1697 245 1703 248
rect 1710 245 1712 249
rect 1716 245 1719 249
rect 1697 241 1698 245
rect 1702 241 1703 245
rect 1715 241 1719 245
rect 1729 244 1735 251
rect 1739 255 1756 256
rect 1743 251 1756 255
rect 1739 250 1756 251
rect 1748 242 1756 250
rect 1697 237 1706 241
rect 1710 237 1711 241
rect 1715 237 1731 241
rect 1735 237 1736 241
rect 1752 238 1756 242
rect 1697 236 1711 237
rect 1698 224 1701 236
rect 1698 221 1741 224
rect 1684 187 1688 191
rect 1684 175 1692 187
rect 1697 211 1701 212
rect 1697 189 1701 207
rect 1705 210 1725 212
rect 1729 210 1742 212
rect 1705 208 1742 210
rect 1705 201 1709 208
rect 1720 203 1721 204
rect 1705 196 1709 197
rect 1713 200 1721 203
rect 1725 203 1726 204
rect 1725 200 1734 203
rect 1713 199 1734 200
rect 1713 192 1717 199
rect 1712 191 1717 192
rect 1697 185 1706 189
rect 1716 187 1717 191
rect 1712 186 1717 187
rect 1721 194 1725 195
rect 1702 182 1706 185
rect 1721 182 1725 190
rect 1702 178 1725 182
rect 1730 183 1734 199
rect 1738 193 1742 208
rect 1738 188 1742 189
rect 1748 211 1756 238
rect 1762 246 1768 249
rect 1762 214 1765 246
rect 1752 207 1756 211
rect 1748 201 1762 207
rect 1779 203 1784 271
rect 1748 197 1758 201
rect 1767 202 1812 203
rect 1767 198 1770 202
rect 1774 199 1806 202
rect 1774 198 1775 199
rect 1805 198 1806 199
rect 1810 198 1812 202
rect 1748 193 1762 197
rect 1748 192 1774 193
rect 1748 188 1770 192
rect 1748 187 1774 188
rect 1777 191 1785 195
rect 1789 191 1804 195
rect 1730 179 1736 183
rect 1740 179 1741 183
rect 1684 171 1691 175
rect 1695 171 1698 175
rect 1702 171 1703 175
rect 1581 140 1586 142
rect 1534 139 1590 140
rect 1538 135 1590 139
rect 1451 105 1457 109
rect 1461 105 1467 109
rect 1471 105 1487 109
rect 1497 106 1498 112
rect 1403 97 1406 102
rect 1424 101 1487 105
rect 1424 97 1429 101
rect 1164 94 1429 97
rect 1581 97 1586 135
rect 1684 109 1692 171
rect 1710 165 1714 178
rect 1748 173 1762 187
rect 1777 182 1781 191
rect 1792 185 1796 188
rect 1769 178 1770 182
rect 1774 178 1781 182
rect 1800 187 1804 191
rect 1808 190 1812 198
rect 1818 201 1826 207
rect 1822 197 1826 201
rect 1818 191 1826 197
rect 1815 190 1826 191
rect 1800 183 1812 187
rect 1819 186 1826 190
rect 1815 185 1826 186
rect 1784 175 1788 180
rect 1792 179 1796 181
rect 1792 175 1805 179
rect 1722 169 1727 173
rect 1731 169 1735 173
rect 1748 172 1758 173
rect 1722 167 1735 169
rect 1697 157 1703 164
rect 1710 161 1712 165
rect 1716 161 1719 165
rect 1729 163 1735 167
rect 1739 171 1758 172
rect 1743 169 1758 171
rect 1762 172 1774 173
rect 1762 169 1770 172
rect 1743 168 1770 169
rect 1743 167 1774 168
rect 1777 171 1780 174
rect 1802 171 1805 175
rect 1781 167 1793 171
rect 1801 167 1805 171
rect 1808 172 1812 183
rect 1808 167 1812 168
rect 1739 166 1762 167
rect 1715 157 1719 161
rect 1729 160 1744 163
rect 1697 153 1706 157
rect 1710 153 1711 157
rect 1715 153 1731 157
rect 1735 153 1736 157
rect 1697 152 1711 153
rect 1707 147 1710 152
rect 1707 144 1724 147
rect 1741 136 1744 160
rect 1748 159 1756 166
rect 1818 163 1826 185
rect 1874 173 1878 274
rect 1874 170 1879 173
rect 1768 159 1777 162
rect 1790 159 1812 162
rect 1823 159 1827 163
rect 1748 158 1761 159
rect 1752 154 1761 158
rect 1774 155 1777 159
rect 1748 144 1761 154
rect 1766 154 1806 155
rect 1766 150 1767 154
rect 1771 151 1795 154
rect 1771 150 1772 151
rect 1794 150 1795 151
rect 1799 150 1802 154
rect 1776 147 1780 148
rect 1748 140 1763 144
rect 1767 140 1768 144
rect 1809 145 1812 159
rect 1684 108 1709 109
rect 1684 104 1688 108
rect 1692 105 1709 108
rect 1713 105 1714 109
rect 1721 106 1724 110
rect 1728 106 1735 110
rect 1730 105 1735 106
rect 1684 94 1692 104
rect 1684 90 1688 94
rect 1684 86 1692 90
rect 1697 98 1698 102
rect 1702 98 1703 102
rect 1734 101 1735 105
rect 1697 96 1703 98
rect 1697 92 1698 96
rect 1702 95 1703 96
rect 1713 99 1726 100
rect 1717 95 1726 99
rect 1730 97 1735 101
rect 1739 108 1743 109
rect 1702 92 1710 95
rect 1713 94 1726 95
rect 1739 94 1743 104
rect 1697 89 1710 92
rect 1722 90 1743 94
rect 1748 90 1761 140
rect 1766 134 1770 135
rect 1776 134 1780 143
rect 1817 144 1827 159
rect 1815 143 1827 144
rect 1785 137 1786 141
rect 1790 138 1803 141
rect 1819 139 1827 143
rect 1815 138 1827 139
rect 1790 137 1807 138
rect 1799 135 1807 137
rect 1766 114 1770 130
rect 1774 130 1795 134
rect 1774 124 1778 130
rect 1791 127 1795 130
rect 1799 127 1800 131
rect 1774 119 1778 120
rect 1782 123 1783 127
rect 1787 124 1788 127
rect 1787 123 1795 124
rect 1782 119 1795 123
rect 1803 119 1807 135
rect 1766 110 1767 114
rect 1771 110 1774 114
rect 1778 110 1779 114
rect 1783 108 1787 112
rect 1767 104 1771 105
rect 1774 104 1783 107
rect 1774 103 1787 104
rect 1767 99 1771 100
rect 1783 101 1787 103
rect 1767 95 1779 99
rect 1713 89 1717 90
rect 1083 83 1478 84
rect 1083 79 1626 83
rect 1684 85 1713 86
rect 1684 82 1717 85
rect 1722 86 1726 90
rect 1752 88 1761 90
rect 1752 87 1764 88
rect 1752 86 1760 87
rect 1655 77 1674 80
rect 1684 80 1692 82
rect 1722 81 1726 82
rect 1684 76 1688 80
rect 1737 79 1743 86
rect 1712 78 1713 79
rect 1338 71 1673 72
rect 1068 69 1674 71
rect 1068 68 1351 69
rect 1356 60 1395 61
rect 1561 60 1650 62
rect 1356 56 1650 60
rect 1655 56 1656 62
rect 992 44 1528 48
rect 1196 43 1528 44
rect 1156 34 1624 35
rect 1063 31 1624 34
rect 1063 30 1342 31
rect 1618 30 1624 31
rect 1063 29 1170 30
rect 1618 29 1621 30
rect 1403 18 1516 22
rect 1403 17 1523 18
rect 1670 3 1674 69
rect 1684 44 1692 76
rect 1705 75 1713 78
rect 1717 78 1718 79
rect 1735 78 1736 79
rect 1717 75 1726 78
rect 1705 74 1726 75
rect 1730 75 1736 78
rect 1740 75 1743 79
rect 1730 74 1743 75
rect 1748 83 1760 86
rect 1748 82 1764 83
rect 1767 87 1771 92
rect 1748 80 1761 82
rect 1752 76 1761 80
rect 1748 73 1761 76
rect 1753 59 1761 73
rect 1767 76 1771 83
rect 1775 83 1779 95
rect 1783 94 1787 97
rect 1791 91 1795 119
rect 1782 87 1783 91
rect 1787 87 1795 91
rect 1791 86 1795 87
rect 1799 115 1807 119
rect 1799 96 1803 115
rect 1817 109 1827 138
rect 1807 108 1827 109
rect 1811 104 1814 108
rect 1818 104 1827 108
rect 1807 103 1827 104
rect 1803 92 1806 96
rect 1810 92 1811 96
rect 1799 83 1803 92
rect 1817 87 1827 103
rect 1775 81 1803 83
rect 1807 86 1827 87
rect 1811 82 1814 86
rect 1818 82 1827 86
rect 1807 81 1827 82
rect 1775 79 1783 81
rect 1782 77 1783 79
rect 1787 79 1803 81
rect 1787 77 1788 79
rect 1791 74 1792 76
rect 1771 72 1792 74
rect 1796 72 1799 76
rect 1803 72 1804 76
rect 1767 70 1804 72
rect 1797 58 1800 70
rect 1817 66 1827 81
rect 1807 63 1827 66
rect 1701 52 1735 56
rect 1799 54 1800 55
rect 1807 54 1810 63
rect 1817 59 1827 63
rect 1799 51 1810 54
rect 1799 50 1800 51
rect 1823 44 1827 59
rect 1684 40 1827 44
rect 1803 39 1827 40
rect 1702 30 1717 34
rect 1740 34 1792 37
rect 1875 35 1879 170
rect 1886 58 1889 329
rect 1921 258 1925 369
rect 1941 368 1956 369
rect 1955 349 1959 356
rect 1955 348 1960 349
rect 1955 344 1956 348
rect 1963 348 1967 369
rect 1970 363 1983 364
rect 1970 359 1973 363
rect 1977 359 1979 363
rect 1970 358 1983 359
rect 1970 351 1976 358
rect 1986 352 1990 369
rect 2056 369 2068 370
rect 2072 370 2152 373
rect 2072 369 2136 370
rect 2033 358 2045 364
rect 2052 363 2056 366
rect 2140 369 2152 370
rect 2156 369 2189 373
rect 2193 369 2203 373
rect 2207 369 2217 373
rect 2221 371 2286 373
rect 2290 371 2300 375
rect 2304 371 2314 375
rect 2318 372 2397 375
rect 2318 371 2381 372
rect 2221 369 2256 371
rect 2066 360 2088 364
rect 2092 360 2093 364
rect 2117 363 2129 364
rect 2066 359 2070 360
rect 2052 358 2056 359
rect 2033 355 2038 358
rect 2033 354 2034 355
rect 1963 344 1966 348
rect 1970 344 1971 348
rect 1975 344 1976 348
rect 1980 344 1981 348
rect 1986 347 1990 348
rect 2025 351 2034 354
rect 2059 355 2070 359
rect 2117 359 2122 363
rect 2126 359 2129 363
rect 2117 358 2129 359
rect 2136 363 2140 366
rect 2150 360 2172 364
rect 2176 360 2177 364
rect 2150 359 2154 360
rect 2136 358 2140 359
rect 2059 351 2063 355
rect 2077 352 2078 356
rect 2082 352 2093 356
rect 1955 343 1960 344
rect 1955 335 1959 343
rect 1975 339 1981 344
rect 1962 335 1963 339
rect 1967 335 1981 339
rect 1987 337 1991 340
rect 2025 337 2028 351
rect 2033 350 2038 351
rect 2042 349 2063 351
rect 1955 326 1959 331
rect 1955 325 1960 326
rect 1955 321 1956 325
rect 1960 321 1967 324
rect 1955 318 1967 321
rect 1971 322 1975 335
rect 2034 345 2042 346
rect 2046 347 2063 349
rect 2034 342 2046 345
rect 1987 331 1991 333
rect 1978 327 1982 331
rect 1986 327 1991 331
rect 1978 326 1991 327
rect 2034 330 2038 342
rect 2059 340 2063 347
rect 2067 345 2068 349
rect 2072 348 2073 349
rect 2072 345 2084 348
rect 2067 344 2084 345
rect 2080 341 2084 344
rect 2080 340 2085 341
rect 2048 334 2054 339
rect 2059 336 2071 340
rect 2075 336 2076 340
rect 2080 336 2081 340
rect 2048 332 2050 334
rect 2041 330 2050 332
rect 2080 335 2085 336
rect 2089 336 2093 352
rect 2117 355 2122 358
rect 2117 351 2118 355
rect 2143 355 2154 359
rect 2143 351 2147 355
rect 2161 352 2162 356
rect 2166 352 2176 356
rect 2117 350 2122 351
rect 2126 349 2147 351
rect 2118 345 2126 346
rect 2130 347 2147 349
rect 2118 342 2130 345
rect 2080 331 2084 335
rect 2041 326 2054 330
rect 2060 327 2084 331
rect 2089 332 2091 336
rect 2034 325 2038 326
rect 2060 325 2064 327
rect 1971 318 1985 322
rect 1989 318 1990 322
rect 2047 318 2048 322
rect 2052 318 2053 322
rect 2089 323 2093 332
rect 2118 330 2122 342
rect 2143 340 2147 347
rect 2151 345 2152 349
rect 2156 348 2157 349
rect 2156 345 2168 348
rect 2151 344 2168 345
rect 2164 341 2168 344
rect 2164 340 2169 341
rect 2132 334 2138 339
rect 2143 336 2155 340
rect 2159 336 2160 340
rect 2164 336 2165 340
rect 2132 332 2134 334
rect 2125 330 2134 332
rect 2164 335 2169 336
rect 2164 331 2168 335
rect 2125 326 2138 330
rect 2144 327 2168 331
rect 2118 325 2122 326
rect 2144 325 2148 327
rect 2060 320 2064 321
rect 2069 319 2070 323
rect 2074 319 2093 323
rect 2047 313 2053 318
rect 2131 318 2132 322
rect 2136 318 2137 322
rect 2173 323 2177 352
rect 2187 349 2191 356
rect 2187 348 2192 349
rect 2187 344 2188 348
rect 2195 348 2199 369
rect 2202 363 2215 364
rect 2202 359 2205 363
rect 2209 359 2211 363
rect 2202 358 2215 359
rect 2202 351 2208 358
rect 2218 352 2222 369
rect 2195 344 2198 348
rect 2202 344 2203 348
rect 2207 344 2208 348
rect 2212 344 2213 348
rect 2218 347 2222 348
rect 2187 343 2192 344
rect 2187 335 2191 343
rect 2207 339 2213 344
rect 2194 335 2195 339
rect 2199 335 2213 339
rect 2219 338 2223 340
rect 2144 320 2148 321
rect 2153 319 2154 323
rect 2158 319 2177 323
rect 2181 332 2191 335
rect 2181 320 2184 332
rect 2131 313 2137 318
rect 2187 326 2191 332
rect 2187 325 2192 326
rect 2187 321 2188 325
rect 2192 321 2199 324
rect 2187 318 2199 321
rect 2203 322 2207 335
rect 2219 331 2223 334
rect 2210 327 2214 331
rect 2218 327 2223 331
rect 2210 326 2223 327
rect 2203 318 2217 322
rect 2221 318 2222 322
rect 1954 309 1957 313
rect 1961 309 1967 313
rect 1971 309 2035 313
rect 2039 309 2088 313
rect 2092 309 2119 313
rect 2123 309 2172 313
rect 2176 309 2189 313
rect 2193 309 2199 313
rect 2203 312 2227 313
rect 2203 309 2221 312
rect 1940 306 2221 309
rect 1940 305 2227 306
rect 2044 303 2088 305
rect 2044 299 2050 303
rect 2054 299 2078 303
rect 2082 299 2088 303
rect 2241 299 2244 361
rect 2048 291 2054 299
rect 2048 287 2049 291
rect 2053 287 2054 291
rect 2059 291 2063 292
rect 2068 291 2074 299
rect 2241 294 2242 299
rect 2068 287 2069 291
rect 2073 287 2074 291
rect 2079 291 2084 294
rect 2083 287 2084 291
rect 2059 284 2063 287
rect 2079 286 2084 287
rect 2059 280 2076 284
rect 2048 268 2052 278
rect 2056 273 2061 277
rect 2072 276 2076 280
rect 2056 265 2062 269
rect 2066 265 2069 269
rect 1920 238 1925 258
rect 2056 259 2060 265
rect 2072 261 2076 272
rect 2043 256 2060 259
rect 2064 257 2076 261
rect 2080 282 2241 286
rect 2064 253 2068 257
rect 2080 256 2084 282
rect 2250 260 2254 369
rect 2284 351 2288 358
rect 2284 350 2289 351
rect 2284 346 2285 350
rect 2292 350 2296 371
rect 2299 365 2312 366
rect 2299 361 2302 365
rect 2306 361 2308 365
rect 2299 360 2312 361
rect 2299 353 2305 360
rect 2315 354 2319 371
rect 2385 371 2397 372
rect 2401 372 2481 375
rect 2401 371 2465 372
rect 2362 360 2374 366
rect 2381 365 2385 368
rect 2469 371 2481 372
rect 2485 371 2518 375
rect 2522 371 2532 375
rect 2536 371 2546 375
rect 2550 374 2613 375
rect 2617 374 2627 378
rect 2631 374 2641 378
rect 2645 375 2724 378
rect 2645 374 2708 375
rect 2550 371 2586 374
rect 2395 362 2417 366
rect 2421 362 2422 366
rect 2437 365 2458 366
rect 2395 361 2399 362
rect 2381 360 2385 361
rect 2362 357 2367 360
rect 2362 356 2363 357
rect 2292 346 2295 350
rect 2299 346 2300 350
rect 2304 346 2305 350
rect 2309 346 2310 350
rect 2315 349 2319 350
rect 2354 353 2363 356
rect 2388 357 2399 361
rect 2437 361 2451 365
rect 2455 361 2458 365
rect 2437 360 2458 361
rect 2465 365 2469 368
rect 2479 362 2501 366
rect 2505 362 2506 366
rect 2479 361 2483 362
rect 2465 360 2469 361
rect 2388 353 2392 357
rect 2406 354 2407 358
rect 2411 354 2422 358
rect 2284 345 2289 346
rect 2284 337 2288 345
rect 2304 341 2310 346
rect 2291 337 2292 341
rect 2296 337 2310 341
rect 2316 339 2320 342
rect 2354 339 2357 353
rect 2362 352 2367 353
rect 2371 351 2392 353
rect 2284 328 2288 333
rect 2284 327 2289 328
rect 2284 323 2285 327
rect 2289 323 2296 326
rect 2284 320 2296 323
rect 2300 324 2304 337
rect 2363 347 2371 348
rect 2375 349 2392 351
rect 2363 344 2375 347
rect 2316 333 2320 335
rect 2307 329 2311 333
rect 2315 329 2320 333
rect 2307 328 2320 329
rect 2363 332 2367 344
rect 2388 342 2392 349
rect 2396 347 2397 351
rect 2401 350 2402 351
rect 2401 347 2413 350
rect 2396 346 2413 347
rect 2409 343 2413 346
rect 2409 342 2414 343
rect 2377 336 2383 341
rect 2388 338 2400 342
rect 2404 338 2405 342
rect 2409 338 2410 342
rect 2377 334 2379 336
rect 2370 332 2379 334
rect 2409 337 2414 338
rect 2418 338 2422 354
rect 2446 357 2451 360
rect 2446 353 2447 357
rect 2472 357 2483 361
rect 2472 353 2476 357
rect 2490 354 2491 358
rect 2495 354 2508 358
rect 2446 352 2451 353
rect 2455 351 2476 353
rect 2447 347 2455 348
rect 2459 349 2476 351
rect 2447 344 2459 347
rect 2409 333 2413 337
rect 2370 328 2383 332
rect 2389 329 2413 333
rect 2418 334 2420 338
rect 2363 327 2367 328
rect 2389 327 2393 329
rect 2300 320 2314 324
rect 2318 320 2319 324
rect 2376 320 2377 324
rect 2381 320 2382 324
rect 2418 325 2422 334
rect 2447 332 2451 344
rect 2472 342 2476 349
rect 2480 347 2481 351
rect 2485 350 2486 351
rect 2485 347 2497 350
rect 2480 346 2497 347
rect 2493 343 2497 346
rect 2493 342 2498 343
rect 2461 336 2467 341
rect 2472 338 2484 342
rect 2488 338 2489 342
rect 2493 338 2494 342
rect 2461 334 2463 336
rect 2454 332 2463 334
rect 2493 337 2498 338
rect 2493 333 2497 337
rect 2454 328 2467 332
rect 2473 329 2497 333
rect 2447 327 2451 328
rect 2473 327 2477 329
rect 2389 322 2393 323
rect 2398 321 2399 325
rect 2403 321 2422 325
rect 2376 315 2382 320
rect 2460 320 2461 324
rect 2465 320 2466 324
rect 2502 325 2506 354
rect 2516 351 2520 358
rect 2516 350 2521 351
rect 2516 346 2517 350
rect 2524 350 2528 371
rect 2531 365 2544 366
rect 2531 361 2534 365
rect 2538 361 2540 365
rect 2531 360 2544 361
rect 2531 353 2537 360
rect 2547 354 2551 371
rect 2524 346 2527 350
rect 2531 346 2532 350
rect 2536 346 2537 350
rect 2541 346 2542 350
rect 2547 349 2551 350
rect 2516 345 2521 346
rect 2516 337 2520 345
rect 2536 341 2542 346
rect 2523 337 2524 341
rect 2528 337 2542 341
rect 2548 340 2552 342
rect 2473 322 2477 323
rect 2482 321 2483 325
rect 2487 321 2506 325
rect 2510 334 2520 337
rect 2510 322 2513 334
rect 2460 315 2466 320
rect 2516 328 2520 334
rect 2516 327 2521 328
rect 2516 323 2517 327
rect 2521 323 2528 326
rect 2516 320 2528 323
rect 2532 324 2536 337
rect 2548 333 2552 336
rect 2539 329 2543 333
rect 2547 329 2552 333
rect 2539 328 2552 329
rect 2532 320 2546 324
rect 2550 320 2551 324
rect 2283 311 2286 315
rect 2290 311 2296 315
rect 2300 311 2364 315
rect 2368 311 2417 315
rect 2421 311 2448 315
rect 2452 311 2501 315
rect 2505 311 2518 315
rect 2522 311 2528 315
rect 2532 314 2556 315
rect 2532 311 2548 314
rect 2283 310 2548 311
rect 2268 308 2548 310
rect 2554 308 2556 314
rect 2268 307 2556 308
rect 2268 306 2284 307
rect 2373 305 2417 307
rect 2373 301 2379 305
rect 2383 301 2407 305
rect 2411 301 2417 305
rect 2079 255 2084 256
rect 2048 249 2049 253
rect 2053 249 2068 253
rect 2071 251 2079 253
rect 2083 251 2084 255
rect 2071 249 2084 251
rect 2066 243 2067 246
rect 2044 242 2067 243
rect 2071 243 2072 246
rect 2071 242 2078 243
rect 2044 239 2078 242
rect 2082 239 2088 243
rect 2044 238 2088 239
rect 2249 240 2254 260
rect 2259 263 2262 294
rect 2377 293 2383 301
rect 2377 289 2378 293
rect 2382 289 2383 293
rect 2388 293 2392 294
rect 2397 293 2403 301
rect 2397 289 2398 293
rect 2402 289 2403 293
rect 2408 293 2413 296
rect 2412 289 2413 293
rect 2388 286 2392 289
rect 2408 288 2413 289
rect 2270 282 2338 286
rect 2388 282 2405 286
rect 2377 270 2381 280
rect 2385 275 2390 279
rect 2401 278 2405 282
rect 2385 267 2391 271
rect 2395 267 2398 271
rect 2259 259 2267 263
rect 2273 259 2274 263
rect 2385 261 2389 267
rect 2401 263 2405 274
rect 2372 258 2389 261
rect 2393 259 2405 263
rect 2409 282 2413 288
rect 2409 279 2560 282
rect 2564 279 2565 282
rect 2393 255 2397 259
rect 2409 258 2413 279
rect 2577 263 2581 371
rect 2611 354 2615 361
rect 2611 353 2616 354
rect 2611 349 2612 353
rect 2619 353 2623 374
rect 2626 368 2639 369
rect 2626 364 2629 368
rect 2633 364 2635 368
rect 2626 363 2639 364
rect 2626 356 2632 363
rect 2642 357 2646 374
rect 2712 374 2724 375
rect 2728 375 2808 378
rect 2728 374 2792 375
rect 2689 363 2701 369
rect 2708 368 2712 371
rect 2796 374 2808 375
rect 2812 374 2845 378
rect 2849 374 2859 378
rect 2863 374 2873 378
rect 2877 374 2883 378
rect 2722 365 2744 369
rect 2748 365 2749 369
rect 2762 368 2785 369
rect 2722 364 2726 365
rect 2762 364 2778 368
rect 2782 364 2785 368
rect 2708 363 2712 364
rect 2689 360 2694 363
rect 2689 359 2690 360
rect 2619 349 2622 353
rect 2626 349 2627 353
rect 2631 349 2632 353
rect 2636 349 2637 353
rect 2642 352 2646 353
rect 2611 348 2616 349
rect 2611 340 2615 348
rect 2631 344 2637 349
rect 2618 340 2619 344
rect 2623 340 2637 344
rect 2643 342 2647 345
rect 2611 331 2615 336
rect 2611 330 2616 331
rect 2611 326 2612 330
rect 2616 326 2623 329
rect 2611 323 2623 326
rect 2627 327 2631 340
rect 2643 336 2647 338
rect 2634 332 2638 336
rect 2642 332 2647 336
rect 2634 331 2647 332
rect 2627 323 2641 327
rect 2645 323 2646 327
rect 2670 325 2674 354
rect 2681 356 2690 359
rect 2715 360 2726 364
rect 2715 356 2719 360
rect 2733 357 2734 361
rect 2738 357 2749 361
rect 2681 342 2684 356
rect 2689 355 2694 356
rect 2698 354 2719 356
rect 2690 350 2698 351
rect 2702 352 2719 354
rect 2690 347 2702 350
rect 2690 335 2694 347
rect 2715 345 2719 352
rect 2723 350 2724 354
rect 2728 353 2729 354
rect 2728 350 2740 353
rect 2723 349 2740 350
rect 2736 346 2740 349
rect 2736 345 2741 346
rect 2704 339 2710 344
rect 2715 341 2727 345
rect 2731 341 2732 345
rect 2736 341 2737 345
rect 2704 337 2706 339
rect 2697 335 2706 337
rect 2736 340 2741 341
rect 2745 341 2749 357
rect 2736 336 2740 340
rect 2697 331 2710 335
rect 2716 332 2740 336
rect 2745 337 2747 341
rect 2690 330 2694 331
rect 2716 330 2720 332
rect 2670 321 2671 325
rect 2703 323 2704 327
rect 2708 323 2709 327
rect 2745 328 2749 337
rect 2716 325 2720 326
rect 2725 324 2726 328
rect 2730 324 2749 328
rect 2756 325 2759 356
rect 2703 318 2709 323
rect 2763 318 2767 364
rect 2773 363 2785 364
rect 2792 368 2796 371
rect 2806 365 2828 369
rect 2832 365 2833 369
rect 2806 364 2810 365
rect 2792 363 2796 364
rect 2773 360 2778 363
rect 2773 356 2774 360
rect 2799 360 2810 364
rect 2799 356 2803 360
rect 2817 357 2818 361
rect 2822 357 2833 361
rect 2773 355 2778 356
rect 2782 354 2803 356
rect 2774 350 2782 351
rect 2786 352 2803 354
rect 2774 347 2786 350
rect 2774 335 2778 347
rect 2799 345 2803 352
rect 2807 350 2808 354
rect 2812 353 2813 354
rect 2812 350 2824 353
rect 2807 349 2824 350
rect 2820 346 2824 349
rect 2820 345 2825 346
rect 2788 339 2794 344
rect 2799 341 2811 345
rect 2815 341 2816 345
rect 2820 341 2821 345
rect 2788 337 2790 339
rect 2781 335 2790 337
rect 2820 340 2825 341
rect 2820 336 2824 340
rect 2781 331 2794 335
rect 2800 332 2824 336
rect 2774 330 2778 331
rect 2800 330 2804 332
rect 2787 323 2788 327
rect 2792 323 2793 327
rect 2829 328 2833 357
rect 2843 354 2847 361
rect 2843 353 2848 354
rect 2843 349 2844 353
rect 2851 353 2855 374
rect 2858 368 2871 369
rect 2858 364 2861 368
rect 2865 364 2867 368
rect 2858 363 2871 364
rect 2858 356 2864 363
rect 2874 357 2878 374
rect 2851 349 2854 353
rect 2858 349 2859 353
rect 2863 349 2864 353
rect 2868 349 2869 353
rect 2874 352 2878 353
rect 2843 348 2848 349
rect 2843 340 2847 348
rect 2863 344 2869 349
rect 2850 340 2851 344
rect 2855 340 2869 344
rect 2875 343 2879 345
rect 2800 325 2804 326
rect 2809 324 2810 328
rect 2814 324 2833 328
rect 2837 337 2847 340
rect 2837 325 2840 337
rect 2787 318 2793 323
rect 2843 331 2847 337
rect 2843 330 2848 331
rect 2843 326 2844 330
rect 2848 326 2855 329
rect 2843 323 2855 326
rect 2859 327 2863 340
rect 2875 336 2879 339
rect 2866 332 2870 336
rect 2874 332 2879 336
rect 2866 331 2879 332
rect 2859 323 2873 327
rect 2877 323 2878 327
rect 2610 317 2613 318
rect 2608 314 2613 317
rect 2617 314 2623 318
rect 2627 314 2691 318
rect 2695 314 2744 318
rect 2748 314 2775 318
rect 2779 314 2828 318
rect 2832 314 2845 318
rect 2849 314 2855 318
rect 2859 314 2883 318
rect 2608 312 2883 314
rect 2595 310 2883 312
rect 2595 309 2612 310
rect 2595 308 2611 309
rect 2700 308 2744 310
rect 2700 304 2706 308
rect 2710 304 2734 308
rect 2738 304 2744 308
rect 2704 296 2710 304
rect 2704 292 2705 296
rect 2709 292 2710 296
rect 2715 296 2719 297
rect 2724 296 2730 304
rect 2724 292 2725 296
rect 2729 292 2730 296
rect 2735 296 2740 299
rect 2739 292 2740 296
rect 2596 279 2663 282
rect 2667 279 2668 282
rect 2408 257 2413 258
rect 2377 251 2378 255
rect 2382 251 2397 255
rect 2400 253 2408 255
rect 2412 253 2413 257
rect 2400 251 2413 253
rect 2395 245 2396 248
rect 2373 244 2396 245
rect 2400 245 2401 248
rect 2400 244 2407 245
rect 2373 241 2407 244
rect 2411 241 2417 245
rect 2373 240 2417 241
rect 1920 235 2088 238
rect 1920 234 2048 235
rect 2226 234 2241 238
rect 2045 231 2048 234
rect 2249 237 2417 240
rect 2576 243 2581 263
rect 2673 251 2677 291
rect 2715 289 2719 292
rect 2735 291 2740 292
rect 2715 285 2732 289
rect 2685 257 2688 284
rect 2704 273 2708 283
rect 2712 278 2717 282
rect 2728 281 2732 285
rect 2712 270 2718 274
rect 2722 270 2725 274
rect 2712 264 2716 270
rect 2728 266 2732 277
rect 2699 261 2716 264
rect 2720 262 2732 266
rect 2736 287 2740 291
rect 2736 284 2748 287
rect 2720 258 2724 262
rect 2736 261 2740 284
rect 2756 263 2759 278
rect 2735 260 2740 261
rect 2704 254 2705 258
rect 2709 254 2724 258
rect 2727 256 2735 258
rect 2739 256 2740 260
rect 2727 254 2740 256
rect 2722 248 2723 251
rect 2673 246 2677 247
rect 2700 247 2723 248
rect 2727 248 2728 251
rect 2755 250 2760 263
rect 2727 247 2734 248
rect 2700 244 2734 247
rect 2738 244 2744 248
rect 2700 243 2744 244
rect 2910 248 2913 401
rect 2870 245 2913 248
rect 2576 240 2744 243
rect 2576 239 2700 240
rect 2249 236 2375 237
rect 2705 236 2708 240
rect 2372 233 2375 236
rect 2576 233 2882 236
rect 1920 227 2226 231
rect 1920 223 1956 227
rect 1960 223 1970 227
rect 1974 223 1984 227
rect 1988 224 2067 227
rect 1988 223 2051 224
rect 1920 112 1924 223
rect 1954 203 1958 210
rect 1954 202 1959 203
rect 1954 198 1955 202
rect 1962 202 1966 223
rect 1969 217 1982 218
rect 1969 213 1972 217
rect 1976 213 1978 217
rect 1969 212 1982 213
rect 1969 205 1975 212
rect 1985 206 1989 223
rect 2055 223 2067 224
rect 2071 224 2151 227
rect 2071 223 2135 224
rect 2032 212 2044 218
rect 2051 217 2055 220
rect 2139 223 2151 224
rect 2155 223 2188 227
rect 2192 223 2202 227
rect 2206 223 2216 227
rect 2220 223 2226 227
rect 2249 229 2555 233
rect 2249 225 2285 229
rect 2289 225 2299 229
rect 2303 225 2313 229
rect 2317 226 2396 229
rect 2317 225 2380 226
rect 2065 214 2087 218
rect 2091 214 2092 218
rect 2116 217 2128 218
rect 2104 214 2121 217
rect 2065 213 2069 214
rect 2051 212 2055 213
rect 2032 209 2037 212
rect 2032 208 2033 209
rect 1962 198 1965 202
rect 1969 198 1970 202
rect 1974 198 1975 202
rect 1979 198 1980 202
rect 1985 201 1989 202
rect 2024 205 2033 208
rect 2058 209 2069 213
rect 2058 205 2062 209
rect 2076 206 2077 210
rect 2081 206 2092 210
rect 1954 197 1959 198
rect 1954 189 1958 197
rect 1974 193 1980 198
rect 1961 189 1962 193
rect 1966 189 1980 193
rect 1986 191 1990 194
rect 2024 191 2027 205
rect 2032 204 2037 205
rect 2041 203 2062 205
rect 1954 180 1958 185
rect 1954 179 1959 180
rect 1954 175 1955 179
rect 1959 175 1966 178
rect 1954 172 1966 175
rect 1970 176 1974 189
rect 2033 199 2041 200
rect 2045 201 2062 203
rect 2033 196 2045 199
rect 1986 185 1990 187
rect 1977 181 1981 185
rect 1985 181 1990 185
rect 1977 180 1990 181
rect 2033 184 2037 196
rect 2058 194 2062 201
rect 2066 199 2067 203
rect 2071 202 2072 203
rect 2071 199 2083 202
rect 2066 198 2083 199
rect 2079 195 2083 198
rect 2079 194 2084 195
rect 2047 188 2053 193
rect 2058 190 2070 194
rect 2074 190 2075 194
rect 2079 190 2080 194
rect 2047 186 2049 188
rect 2040 184 2049 186
rect 2079 189 2084 190
rect 2088 190 2092 206
rect 2079 185 2083 189
rect 2040 180 2053 184
rect 2059 181 2083 185
rect 2088 186 2090 190
rect 2033 179 2037 180
rect 2059 179 2063 181
rect 1970 172 1984 176
rect 1988 172 1989 176
rect 2046 172 2047 176
rect 2051 172 2052 176
rect 2088 177 2092 186
rect 2059 174 2063 175
rect 2068 173 2069 177
rect 2073 173 2092 177
rect 2104 174 2107 214
rect 2116 213 2121 214
rect 2125 213 2128 217
rect 2116 212 2128 213
rect 2135 217 2139 220
rect 2149 214 2171 218
rect 2175 214 2176 218
rect 2149 213 2153 214
rect 2135 212 2139 213
rect 2116 209 2121 212
rect 2116 205 2117 209
rect 2142 209 2153 213
rect 2142 205 2146 209
rect 2160 206 2161 210
rect 2165 206 2176 210
rect 2116 204 2121 205
rect 2125 203 2146 205
rect 2117 199 2125 200
rect 2129 201 2146 203
rect 2117 196 2129 199
rect 2117 184 2121 196
rect 2142 194 2146 201
rect 2150 199 2151 203
rect 2155 202 2156 203
rect 2155 199 2167 202
rect 2150 198 2167 199
rect 2163 195 2167 198
rect 2172 197 2176 206
rect 2186 203 2190 210
rect 2186 202 2191 203
rect 2186 198 2187 202
rect 2194 202 2198 223
rect 2201 217 2214 218
rect 2201 213 2204 217
rect 2208 213 2210 217
rect 2201 212 2214 213
rect 2201 205 2207 212
rect 2217 206 2221 223
rect 2194 198 2197 202
rect 2201 198 2202 202
rect 2206 198 2207 202
rect 2211 198 2212 202
rect 2217 201 2221 202
rect 2163 194 2168 195
rect 2131 188 2137 193
rect 2142 190 2154 194
rect 2158 190 2159 194
rect 2163 190 2164 194
rect 2131 186 2133 188
rect 2124 184 2133 186
rect 2163 189 2168 190
rect 2172 194 2179 197
rect 2186 197 2191 198
rect 2163 185 2167 189
rect 2124 180 2137 184
rect 2143 181 2167 185
rect 2117 179 2121 180
rect 2143 179 2147 181
rect 2046 167 2052 172
rect 2130 172 2131 176
rect 2135 172 2136 176
rect 2172 177 2176 194
rect 2186 189 2190 197
rect 2206 193 2212 198
rect 2193 189 2194 193
rect 2198 189 2212 193
rect 2218 192 2222 194
rect 2143 174 2147 175
rect 2152 173 2153 177
rect 2157 173 2176 177
rect 2180 186 2190 189
rect 2180 174 2183 186
rect 2130 167 2136 172
rect 2186 180 2190 186
rect 2186 179 2191 180
rect 2186 175 2187 179
rect 2191 175 2198 178
rect 2186 172 2198 175
rect 2202 176 2206 189
rect 2218 185 2222 188
rect 2209 181 2213 185
rect 2217 181 2222 185
rect 2209 180 2222 181
rect 2202 172 2216 176
rect 2220 172 2221 176
rect 1953 163 1956 167
rect 1960 163 1966 167
rect 1970 163 2034 167
rect 2038 163 2087 167
rect 2091 163 2118 167
rect 2122 163 2171 167
rect 2175 163 2188 167
rect 2192 163 2198 167
rect 2202 163 2221 167
rect 1953 160 2221 163
rect 1953 159 2226 160
rect 2043 157 2087 159
rect 2043 153 2049 157
rect 2053 153 2077 157
rect 2081 153 2087 157
rect 2047 145 2053 153
rect 2047 141 2048 145
rect 2052 141 2053 145
rect 2058 145 2062 146
rect 2067 145 2073 153
rect 2174 150 2215 153
rect 2067 141 2068 145
rect 2072 141 2073 145
rect 2078 145 2083 148
rect 2082 141 2083 145
rect 2058 138 2062 141
rect 2078 140 2083 141
rect 2058 134 2075 138
rect 2047 122 2051 132
rect 2055 127 2060 131
rect 2071 130 2075 134
rect 2055 119 2061 123
rect 2065 119 2068 123
rect 1919 92 1924 112
rect 2055 113 2059 119
rect 2071 115 2075 126
rect 2042 110 2059 113
rect 2063 111 2075 115
rect 2079 127 2083 140
rect 2171 132 2194 135
rect 2199 132 2200 135
rect 2079 124 2120 127
rect 2063 107 2067 111
rect 2079 110 2083 124
rect 2078 109 2083 110
rect 2047 103 2048 107
rect 2052 103 2067 107
rect 2070 105 2078 107
rect 2082 105 2083 109
rect 2070 103 2083 105
rect 2065 97 2066 100
rect 2043 96 2066 97
rect 2070 97 2071 100
rect 2070 96 2077 97
rect 2043 93 2077 96
rect 2081 93 2087 97
rect 2043 92 2087 93
rect 1919 89 2087 92
rect 1919 88 2043 89
rect 1967 77 1971 88
rect 2115 83 2119 124
rect 1970 72 1971 77
rect 2113 71 2119 83
rect 1886 57 1908 58
rect 2113 57 2117 71
rect 1886 55 2118 57
rect 1905 53 2118 55
rect 2212 49 2215 150
rect 2224 131 2240 135
rect 2249 114 2253 225
rect 2283 205 2287 212
rect 2283 204 2288 205
rect 2283 200 2284 204
rect 2291 204 2295 225
rect 2298 219 2311 220
rect 2298 215 2301 219
rect 2305 215 2307 219
rect 2298 214 2311 215
rect 2298 207 2304 214
rect 2314 208 2318 225
rect 2384 225 2396 226
rect 2400 226 2480 229
rect 2400 225 2464 226
rect 2361 214 2373 220
rect 2380 219 2384 222
rect 2468 225 2480 226
rect 2484 225 2517 229
rect 2521 225 2531 229
rect 2535 225 2545 229
rect 2549 225 2555 229
rect 2576 232 2832 233
rect 2576 228 2612 232
rect 2616 228 2626 232
rect 2630 228 2640 232
rect 2644 229 2723 232
rect 2644 228 2707 229
rect 2394 216 2416 220
rect 2420 216 2421 220
rect 2445 219 2457 220
rect 2394 215 2398 216
rect 2380 214 2384 215
rect 2361 211 2366 214
rect 2361 210 2362 211
rect 2291 200 2294 204
rect 2298 200 2299 204
rect 2303 200 2304 204
rect 2308 200 2309 204
rect 2314 203 2318 204
rect 2353 207 2362 210
rect 2387 211 2398 215
rect 2445 215 2450 219
rect 2454 215 2457 219
rect 2445 214 2457 215
rect 2464 219 2468 222
rect 2478 216 2500 220
rect 2504 216 2505 220
rect 2478 215 2482 216
rect 2464 214 2468 215
rect 2387 207 2391 211
rect 2405 208 2406 212
rect 2410 208 2421 212
rect 2283 199 2288 200
rect 2283 191 2287 199
rect 2303 195 2309 200
rect 2290 191 2291 195
rect 2295 191 2309 195
rect 2315 193 2319 196
rect 2283 182 2287 187
rect 2283 181 2288 182
rect 2283 177 2284 181
rect 2288 177 2295 180
rect 2283 174 2295 177
rect 2299 178 2303 191
rect 2315 187 2319 189
rect 2306 183 2310 187
rect 2314 183 2319 187
rect 2306 182 2319 183
rect 2299 174 2313 178
rect 2317 174 2318 178
rect 2343 176 2346 196
rect 2353 193 2356 207
rect 2361 206 2366 207
rect 2370 205 2391 207
rect 2362 201 2370 202
rect 2374 203 2391 205
rect 2362 198 2374 201
rect 2362 186 2366 198
rect 2387 196 2391 203
rect 2395 201 2396 205
rect 2400 204 2401 205
rect 2400 201 2412 204
rect 2395 200 2412 201
rect 2408 197 2412 200
rect 2408 196 2413 197
rect 2376 190 2382 195
rect 2387 192 2399 196
rect 2403 192 2404 196
rect 2408 192 2409 196
rect 2376 188 2378 190
rect 2369 186 2378 188
rect 2408 191 2413 192
rect 2417 192 2421 208
rect 2445 211 2450 214
rect 2445 207 2446 211
rect 2471 211 2482 215
rect 2471 207 2475 211
rect 2489 208 2490 212
rect 2494 208 2505 212
rect 2445 206 2450 207
rect 2454 205 2475 207
rect 2446 201 2454 202
rect 2458 203 2475 205
rect 2446 198 2458 201
rect 2408 187 2412 191
rect 2369 182 2382 186
rect 2388 183 2412 187
rect 2417 188 2419 192
rect 2362 181 2366 182
rect 2388 181 2392 183
rect 2375 174 2376 178
rect 2380 174 2381 178
rect 2417 179 2421 188
rect 2446 186 2450 198
rect 2471 196 2475 203
rect 2479 201 2480 205
rect 2484 204 2485 205
rect 2484 201 2496 204
rect 2479 200 2496 201
rect 2492 197 2496 200
rect 2501 199 2505 208
rect 2515 205 2519 212
rect 2515 204 2520 205
rect 2515 200 2516 204
rect 2523 204 2527 225
rect 2530 219 2543 220
rect 2530 215 2533 219
rect 2537 215 2539 219
rect 2530 214 2543 215
rect 2530 207 2536 214
rect 2546 208 2550 225
rect 2523 200 2526 204
rect 2530 200 2531 204
rect 2535 200 2536 204
rect 2540 200 2541 204
rect 2546 203 2550 204
rect 2515 199 2520 200
rect 2492 196 2497 197
rect 2460 190 2466 195
rect 2471 192 2483 196
rect 2487 192 2488 196
rect 2492 192 2493 196
rect 2460 188 2462 190
rect 2453 186 2462 188
rect 2492 191 2497 192
rect 2501 195 2508 199
rect 2492 187 2496 191
rect 2453 182 2466 186
rect 2472 183 2496 187
rect 2446 181 2450 182
rect 2472 181 2476 183
rect 2388 176 2392 177
rect 2397 175 2398 179
rect 2402 175 2421 179
rect 2375 169 2381 174
rect 2459 174 2460 178
rect 2464 174 2465 178
rect 2501 179 2505 195
rect 2515 191 2519 199
rect 2535 195 2541 200
rect 2522 191 2523 195
rect 2527 191 2541 195
rect 2547 194 2551 196
rect 2472 176 2476 177
rect 2481 175 2482 179
rect 2486 175 2505 179
rect 2509 188 2519 191
rect 2509 176 2512 188
rect 2459 169 2465 174
rect 2515 182 2519 188
rect 2515 181 2520 182
rect 2515 177 2516 181
rect 2520 177 2527 180
rect 2515 174 2527 177
rect 2531 178 2535 191
rect 2547 187 2551 190
rect 2538 183 2542 187
rect 2546 183 2551 187
rect 2538 182 2551 183
rect 2531 174 2545 178
rect 2549 174 2550 178
rect 2282 165 2285 169
rect 2289 165 2295 169
rect 2299 165 2363 169
rect 2367 165 2416 169
rect 2420 165 2447 169
rect 2451 165 2500 169
rect 2504 165 2517 169
rect 2521 165 2527 169
rect 2531 165 2555 169
rect 2263 162 2548 165
rect 2282 161 2548 162
rect 2552 161 2555 165
rect 2372 159 2416 161
rect 2372 155 2378 159
rect 2382 155 2406 159
rect 2410 155 2416 159
rect 2343 150 2346 152
rect 2376 147 2382 155
rect 2343 132 2346 146
rect 2376 143 2377 147
rect 2381 143 2382 147
rect 2387 147 2391 148
rect 2396 147 2402 155
rect 2396 143 2397 147
rect 2401 143 2402 147
rect 2407 147 2412 150
rect 2411 143 2412 147
rect 2387 140 2391 143
rect 2407 142 2412 143
rect 2387 136 2404 140
rect 2248 94 2253 114
rect 2315 128 2343 131
rect 2315 102 2319 128
rect 2376 124 2380 134
rect 2384 129 2389 133
rect 2400 132 2404 136
rect 2384 121 2390 125
rect 2394 121 2397 125
rect 2384 115 2388 121
rect 2400 117 2404 128
rect 2371 112 2388 115
rect 2392 113 2404 117
rect 2392 109 2396 113
rect 2408 112 2412 142
rect 2439 138 2521 143
rect 2576 117 2580 228
rect 2610 208 2614 215
rect 2610 207 2615 208
rect 2610 203 2611 207
rect 2618 207 2622 228
rect 2625 222 2638 223
rect 2625 218 2628 222
rect 2632 218 2634 222
rect 2625 217 2638 218
rect 2625 210 2631 217
rect 2641 211 2645 228
rect 2711 228 2723 229
rect 2727 229 2807 232
rect 2727 228 2791 229
rect 2688 217 2700 223
rect 2707 222 2711 225
rect 2795 228 2807 229
rect 2811 228 2832 232
rect 2842 232 2882 233
rect 2721 219 2743 223
rect 2747 219 2748 223
rect 2772 222 2784 223
rect 2721 218 2725 219
rect 2707 217 2711 218
rect 2688 214 2693 217
rect 2688 213 2689 214
rect 2618 203 2621 207
rect 2625 203 2626 207
rect 2630 203 2631 207
rect 2635 203 2636 207
rect 2641 206 2645 207
rect 2680 210 2689 213
rect 2714 214 2725 218
rect 2772 218 2777 222
rect 2781 218 2784 222
rect 2772 217 2784 218
rect 2791 222 2795 225
rect 2842 228 2844 232
rect 2848 228 2858 232
rect 2862 228 2872 232
rect 2876 228 2882 232
rect 2805 219 2827 223
rect 2831 219 2832 223
rect 2805 218 2809 219
rect 2791 217 2795 218
rect 2714 210 2718 214
rect 2732 211 2733 215
rect 2737 211 2748 215
rect 2610 202 2615 203
rect 2610 194 2614 202
rect 2630 198 2636 203
rect 2617 194 2618 198
rect 2622 194 2636 198
rect 2642 196 2646 199
rect 2680 196 2683 210
rect 2688 209 2693 210
rect 2697 208 2718 210
rect 2610 185 2614 190
rect 2610 184 2615 185
rect 2610 180 2611 184
rect 2615 180 2622 183
rect 2610 177 2622 180
rect 2626 181 2630 194
rect 2689 204 2697 205
rect 2701 206 2718 208
rect 2689 201 2701 204
rect 2642 190 2646 192
rect 2633 186 2637 190
rect 2641 186 2646 190
rect 2633 185 2646 186
rect 2689 189 2693 201
rect 2714 199 2718 206
rect 2722 204 2723 208
rect 2727 207 2728 208
rect 2727 204 2739 207
rect 2722 203 2739 204
rect 2735 200 2739 203
rect 2735 199 2740 200
rect 2703 193 2709 198
rect 2714 195 2726 199
rect 2730 195 2731 199
rect 2735 195 2736 199
rect 2703 191 2705 193
rect 2689 184 2693 185
rect 2696 189 2705 191
rect 2735 194 2740 195
rect 2744 195 2748 211
rect 2772 214 2777 217
rect 2772 210 2773 214
rect 2798 214 2809 218
rect 2798 210 2802 214
rect 2816 211 2817 215
rect 2821 211 2832 215
rect 2772 209 2777 210
rect 2781 208 2802 210
rect 2773 204 2781 205
rect 2785 206 2802 208
rect 2773 201 2785 204
rect 2735 190 2739 194
rect 2696 185 2709 189
rect 2715 186 2739 190
rect 2744 191 2746 195
rect 2626 177 2640 181
rect 2644 177 2645 181
rect 2696 180 2699 185
rect 2715 184 2719 186
rect 2685 176 2699 180
rect 2702 177 2703 181
rect 2707 177 2708 181
rect 2744 182 2748 191
rect 2773 189 2777 201
rect 2798 199 2802 206
rect 2806 204 2807 208
rect 2811 207 2812 208
rect 2811 204 2823 207
rect 2806 203 2823 204
rect 2819 200 2823 203
rect 2828 201 2832 211
rect 2835 202 2838 226
rect 2842 208 2846 215
rect 2842 207 2847 208
rect 2842 203 2843 207
rect 2850 207 2854 228
rect 2857 222 2870 223
rect 2857 218 2860 222
rect 2864 218 2866 222
rect 2857 217 2870 218
rect 2857 210 2863 217
rect 2873 211 2877 228
rect 2850 203 2853 207
rect 2857 203 2858 207
rect 2862 203 2863 207
rect 2867 203 2868 207
rect 2873 206 2877 207
rect 2842 202 2847 203
rect 2819 199 2824 200
rect 2787 193 2793 198
rect 2798 195 2810 199
rect 2814 195 2815 199
rect 2819 195 2820 199
rect 2787 191 2789 193
rect 2780 189 2789 191
rect 2819 194 2824 195
rect 2828 198 2835 201
rect 2819 190 2823 194
rect 2780 185 2793 189
rect 2799 186 2823 190
rect 2773 184 2777 185
rect 2799 184 2803 186
rect 2715 179 2719 180
rect 2724 178 2725 182
rect 2729 178 2748 182
rect 2685 172 2689 176
rect 2702 172 2708 177
rect 2786 177 2787 181
rect 2791 177 2792 181
rect 2828 182 2832 198
rect 2842 194 2846 202
rect 2862 198 2868 203
rect 2849 194 2850 198
rect 2854 194 2868 198
rect 2874 197 2878 199
rect 2799 179 2803 180
rect 2808 178 2809 182
rect 2813 178 2832 182
rect 2836 191 2846 194
rect 2836 179 2839 191
rect 2786 172 2792 177
rect 2842 185 2846 191
rect 2842 184 2847 185
rect 2842 180 2843 184
rect 2847 180 2854 183
rect 2842 177 2854 180
rect 2858 181 2862 194
rect 2874 190 2878 193
rect 2865 186 2869 190
rect 2873 186 2878 190
rect 2865 185 2878 186
rect 2858 177 2872 181
rect 2876 177 2877 181
rect 2609 169 2612 172
rect 2608 168 2612 169
rect 2616 168 2622 172
rect 2626 168 2690 172
rect 2694 168 2743 172
rect 2747 168 2774 172
rect 2778 168 2827 172
rect 2831 168 2844 172
rect 2848 168 2854 172
rect 2858 168 2882 172
rect 2608 166 2882 168
rect 2589 165 2882 166
rect 2592 164 2882 165
rect 2592 163 2611 164
rect 2699 162 2743 164
rect 2699 158 2705 162
rect 2709 158 2733 162
rect 2737 158 2743 162
rect 2646 156 2650 157
rect 2590 138 2619 143
rect 2407 111 2412 112
rect 2376 105 2377 109
rect 2381 105 2396 109
rect 2399 107 2407 109
rect 2411 109 2412 111
rect 2411 107 2416 109
rect 2399 105 2416 107
rect 2394 99 2395 102
rect 2372 98 2395 99
rect 2399 99 2400 102
rect 2399 98 2406 99
rect 2372 95 2406 98
rect 2410 95 2416 99
rect 2372 94 2416 95
rect 2248 91 2416 94
rect 2575 97 2580 117
rect 2646 115 2650 152
rect 2703 150 2709 158
rect 2703 146 2704 150
rect 2708 146 2709 150
rect 2714 150 2718 151
rect 2723 150 2729 158
rect 2723 146 2724 150
rect 2728 146 2729 150
rect 2734 150 2739 153
rect 2738 146 2739 150
rect 2714 143 2718 146
rect 2734 145 2739 146
rect 2714 139 2731 143
rect 2703 127 2707 137
rect 2711 132 2716 136
rect 2727 135 2731 139
rect 2711 124 2717 128
rect 2721 124 2724 128
rect 2711 118 2715 124
rect 2727 120 2731 131
rect 2698 115 2715 118
rect 2719 116 2731 120
rect 2735 140 2751 145
rect 2719 112 2723 116
rect 2735 115 2739 140
rect 2734 114 2739 115
rect 2703 108 2704 112
rect 2708 108 2723 112
rect 2726 110 2734 112
rect 2738 110 2739 114
rect 2726 108 2739 110
rect 2721 102 2722 105
rect 2699 101 2722 102
rect 2726 102 2727 105
rect 2726 101 2733 102
rect 2699 98 2733 101
rect 2737 98 2743 102
rect 2699 97 2743 98
rect 2575 94 2743 97
rect 2575 93 2699 94
rect 2248 90 2372 91
rect 2361 83 2365 90
rect 2244 81 2288 83
rect 2337 81 2381 83
rect 2424 81 2468 83
rect 2244 79 2468 81
rect 2244 75 2250 79
rect 2254 78 2343 79
rect 2254 75 2288 78
rect 2337 75 2343 78
rect 2347 78 2430 79
rect 2347 75 2381 78
rect 2424 75 2430 78
rect 2434 75 2468 79
rect 2258 67 2264 75
rect 2258 63 2259 67
rect 2263 63 2264 67
rect 2269 69 2273 70
rect 2278 69 2284 75
rect 2319 69 2330 72
rect 2278 65 2279 69
rect 2283 65 2284 69
rect 2248 62 2253 63
rect 2248 58 2249 62
rect 2269 62 2273 65
rect 2248 55 2253 58
rect 2248 51 2249 55
rect 2248 50 2253 51
rect 2256 58 2269 60
rect 2256 56 2273 58
rect 2280 58 2311 62
rect 2248 49 2252 50
rect 2212 45 2252 49
rect 1799 34 1879 35
rect 1688 18 1747 22
rect 1706 3 1710 8
rect 1742 9 1747 18
rect 1774 15 1777 26
rect 1788 22 1792 34
rect 1802 31 1879 34
rect 2248 32 2252 45
rect 2256 45 2260 56
rect 2271 49 2276 53
rect 2280 49 2284 58
rect 2263 41 2266 45
rect 2270 41 2277 45
rect 2256 37 2260 41
rect 2256 33 2268 37
rect 2272 36 2277 41
rect 2248 31 2253 32
rect 2248 27 2249 31
rect 2253 27 2260 30
rect 2248 24 2260 27
rect 2264 29 2268 33
rect 2271 32 2287 36
rect 2264 25 2279 29
rect 2283 25 2284 29
rect 2307 25 2311 58
rect 2327 59 2330 69
rect 2351 67 2357 75
rect 2351 63 2352 67
rect 2356 63 2357 67
rect 2362 69 2366 70
rect 2371 69 2377 75
rect 2371 65 2372 69
rect 2376 65 2377 69
rect 2438 67 2444 75
rect 2417 66 2433 67
rect 2341 62 2346 63
rect 2341 59 2342 62
rect 2327 58 2342 59
rect 2362 62 2366 65
rect 2327 56 2346 58
rect 1788 19 1837 22
rect 2341 55 2346 56
rect 2341 51 2342 55
rect 2341 50 2346 51
rect 2349 58 2362 60
rect 2349 56 2366 58
rect 2341 32 2345 50
rect 2349 45 2353 56
rect 2373 53 2377 62
rect 2421 62 2433 66
rect 2438 63 2439 67
rect 2443 63 2444 67
rect 2449 69 2453 70
rect 2458 69 2464 75
rect 2458 65 2459 69
rect 2463 65 2464 69
rect 2421 61 2429 62
rect 2428 58 2429 61
rect 2449 62 2453 65
rect 2428 55 2433 58
rect 2364 49 2369 53
rect 2373 49 2384 53
rect 2428 51 2429 55
rect 2428 50 2433 51
rect 2436 58 2449 60
rect 2436 56 2453 58
rect 2356 41 2359 45
rect 2363 41 2370 45
rect 2349 37 2353 41
rect 2349 33 2361 37
rect 2341 31 2346 32
rect 2341 27 2342 31
rect 2346 27 2353 30
rect 2341 24 2353 27
rect 2357 29 2361 33
rect 2365 36 2370 41
rect 2365 32 2380 36
rect 2428 32 2432 50
rect 2436 45 2440 56
rect 2460 53 2464 62
rect 2451 49 2456 53
rect 2460 49 2473 53
rect 2443 41 2446 45
rect 2450 41 2457 45
rect 2436 37 2440 41
rect 2436 33 2448 37
rect 2428 31 2433 32
rect 2357 25 2372 29
rect 2376 25 2377 29
rect 2428 27 2429 31
rect 2433 27 2440 30
rect 2428 24 2440 27
rect 2444 29 2448 33
rect 2452 35 2457 41
rect 2452 32 2465 35
rect 2444 25 2459 29
rect 2463 25 2464 29
rect 1761 12 1812 15
rect 2244 15 2250 19
rect 2254 15 2260 19
rect 2264 15 2288 19
rect 2337 15 2343 19
rect 2347 15 2353 19
rect 2357 15 2381 19
rect 2238 14 2381 15
rect 2424 15 2430 19
rect 2434 15 2440 19
rect 2444 15 2468 19
rect 2424 14 2468 15
rect 2238 12 2468 14
rect 2244 11 2288 12
rect 2337 11 2468 12
rect 1742 3 1849 9
rect 1670 0 1710 3
rect 1878 -3 2103 -1
rect 1884 -5 2103 -3
rect 1884 -8 2298 -5
rect 2099 -9 2300 -8
<< metal2 >>
rect 1500 1121 1506 1122
rect 1499 1120 1602 1121
rect 1883 1120 1887 1121
rect 1499 1116 1887 1120
rect 542 1064 893 1065
rect 1500 1064 1506 1116
rect 1598 1115 1887 1116
rect 1813 1110 1818 1111
rect 1817 1105 1818 1110
rect 1549 1077 1554 1101
rect 1813 1095 1818 1105
rect 1814 1085 1818 1095
rect 1815 1081 1818 1085
rect 542 1060 1506 1064
rect 406 1039 511 1040
rect 406 1037 506 1039
rect 124 1032 153 1036
rect 60 1028 127 1032
rect 60 886 65 1028
rect 134 1021 387 1025
rect 75 963 79 1014
rect 134 986 139 1021
rect 382 1017 386 1021
rect 152 1008 153 1011
rect 157 1008 241 1011
rect 245 1008 334 1011
rect 338 1008 359 1011
rect 356 1005 359 1008
rect 406 1005 410 1037
rect 510 1037 511 1039
rect 456 1025 459 1026
rect 456 1022 505 1025
rect 456 1006 459 1022
rect 517 1007 521 1041
rect 542 1025 547 1060
rect 889 1059 1506 1060
rect 1500 1058 1506 1059
rect 988 1034 989 1039
rect 546 1021 547 1025
rect 559 1022 807 1026
rect 559 1018 563 1022
rect 616 1010 705 1013
rect 614 1009 705 1010
rect 709 1009 792 1013
rect 356 1001 410 1005
rect 238 990 382 993
rect 564 992 711 995
rect 133 982 145 986
rect 238 986 241 990
rect 708 988 711 992
rect 150 982 161 986
rect 290 981 291 984
rect 74 961 79 963
rect 74 925 78 961
rect 218 960 266 963
rect 218 959 275 960
rect 263 956 275 959
rect 288 950 291 981
rect 331 976 334 982
rect 612 984 616 987
rect 331 973 382 976
rect 612 976 615 984
rect 564 973 615 976
rect 708 984 709 988
rect 726 986 745 990
rect 803 988 807 1022
rect 988 998 992 1034
rect 1046 1025 1068 1028
rect 1024 998 1027 1021
rect 1133 1008 1213 1011
rect 1133 1002 1136 1008
rect 1094 999 1136 1002
rect 1209 1002 1212 1008
rect 1233 1006 1292 1009
rect 1024 995 1039 998
rect 1166 998 1187 1001
rect 789 984 797 988
rect 802 986 807 988
rect 802 984 1029 986
rect 609 965 612 973
rect 536 962 547 964
rect 609 962 623 965
rect 536 961 541 962
rect 317 958 541 961
rect 545 958 547 962
rect 317 957 547 958
rect 647 956 650 983
rect 709 974 712 984
rect 803 983 1029 984
rect 816 982 1029 983
rect 1015 974 1019 975
rect 709 970 1019 974
rect 662 962 721 965
rect 552 953 650 956
rect 749 962 1011 965
rect 735 958 739 961
rect 735 955 802 958
rect 240 949 293 950
rect 158 946 293 949
rect 552 948 556 953
rect 158 940 161 946
rect 107 937 172 940
rect 74 921 115 925
rect 111 914 115 921
rect 64 882 65 886
rect 72 912 75 913
rect 72 909 79 912
rect 72 844 75 909
rect 115 910 148 913
rect 168 913 171 937
rect 250 937 335 940
rect 339 937 361 940
rect 436 939 501 942
rect 308 927 350 930
rect 358 920 361 937
rect 497 936 501 939
rect 552 936 555 948
rect 798 945 802 955
rect 559 942 579 944
rect 559 941 575 942
rect 559 937 560 941
rect 564 938 575 941
rect 579 939 664 942
rect 763 942 828 945
rect 564 937 579 938
rect 559 936 567 937
rect 394 930 461 933
rect 369 927 397 930
rect 497 933 555 936
rect 357 916 361 920
rect 219 909 252 912
rect 232 905 235 909
rect 344 905 347 911
rect 232 902 347 905
rect 308 893 309 896
rect 306 845 309 893
rect 357 887 360 916
rect 401 911 408 914
rect 351 883 385 887
rect 345 882 385 883
rect 72 841 166 844
rect 176 842 319 845
rect 163 837 166 841
rect 314 811 345 815
rect 295 810 319 811
rect 252 807 319 810
rect 252 806 255 807
rect 196 803 255 806
rect 196 794 200 803
rect 358 796 361 882
rect 369 859 390 863
rect 401 846 404 911
rect 444 912 477 915
rect 497 915 500 933
rect 636 931 794 934
rect 452 898 453 903
rect 452 855 455 898
rect 462 863 466 912
rect 548 911 581 914
rect 561 907 564 911
rect 673 907 676 913
rect 561 904 676 907
rect 728 914 735 917
rect 637 895 638 898
rect 552 874 555 875
rect 552 871 622 874
rect 552 862 555 871
rect 500 859 555 862
rect 500 855 503 859
rect 452 852 504 855
rect 635 847 638 895
rect 678 885 712 889
rect 672 884 712 885
rect 688 856 716 859
rect 728 849 731 914
rect 771 915 804 918
rect 824 918 827 942
rect 906 942 991 945
rect 883 934 957 936
rect 883 933 961 934
rect 787 860 791 915
rect 875 914 908 917
rect 888 910 891 914
rect 1000 910 1003 916
rect 888 907 1003 910
rect 796 873 799 898
rect 964 898 965 901
rect 813 861 872 864
rect 880 860 884 898
rect 962 850 965 898
rect 401 843 495 846
rect 505 844 648 847
rect 728 846 822 849
rect 832 847 975 850
rect 492 839 495 843
rect 819 842 822 846
rect 790 835 810 838
rect 790 833 793 835
rect 550 830 793 833
rect 807 834 810 835
rect 870 835 918 838
rect 807 830 809 834
rect 813 830 814 833
rect 550 814 553 830
rect 870 826 873 835
rect 801 824 873 826
rect 797 823 873 824
rect 879 817 884 820
rect 370 811 553 814
rect 579 813 884 817
rect 579 812 702 813
rect 580 796 585 812
rect 912 799 915 835
rect 106 791 200 794
rect 71 763 78 766
rect 71 698 74 763
rect 114 764 147 767
rect 167 767 170 791
rect 249 791 334 794
rect 358 793 362 796
rect 304 782 351 785
rect 304 775 307 782
rect 359 776 362 793
rect 435 793 500 796
rect 358 773 362 776
rect 467 777 470 793
rect 128 729 131 764
rect 218 763 251 766
rect 231 759 234 763
rect 343 759 346 765
rect 231 756 346 759
rect 307 747 308 750
rect 228 731 231 747
rect 128 725 221 729
rect 227 728 294 731
rect 216 712 221 725
rect 216 708 289 712
rect 305 699 308 747
rect 358 743 361 773
rect 400 765 407 768
rect 353 742 383 743
rect 353 737 382 742
rect 323 708 343 712
rect 71 695 165 698
rect 175 696 318 699
rect 162 691 165 695
rect 224 584 225 588
rect 354 594 360 737
rect 368 728 391 731
rect 381 712 385 713
rect 369 708 385 712
rect 381 687 385 708
rect 400 700 403 765
rect 443 766 476 769
rect 496 769 499 793
rect 578 793 663 796
rect 762 796 827 799
rect 711 788 722 789
rect 633 785 722 788
rect 633 781 636 785
rect 458 719 461 766
rect 547 765 580 768
rect 560 761 563 765
rect 672 761 675 767
rect 560 758 675 761
rect 718 755 721 785
rect 727 768 734 771
rect 467 753 470 754
rect 636 749 637 752
rect 717 751 723 755
rect 467 727 470 749
rect 458 715 557 719
rect 634 701 637 749
rect 676 739 712 742
rect 650 715 709 720
rect 400 697 494 700
rect 504 698 647 701
rect 491 693 494 697
rect 381 683 458 687
rect 455 679 458 683
rect 538 682 540 687
rect 538 679 543 682
rect 413 675 426 678
rect 413 665 416 675
rect 413 662 428 665
rect 439 650 443 675
rect 455 675 543 679
rect 455 674 458 675
rect 454 661 628 664
rect 720 659 723 751
rect 727 703 730 768
rect 770 769 803 772
rect 823 772 826 796
rect 905 796 990 799
rect 998 790 1001 820
rect 968 787 1001 790
rect 968 782 972 787
rect 963 779 972 782
rect 790 733 794 769
rect 874 768 907 771
rect 887 764 890 768
rect 999 764 1002 770
rect 887 761 1002 764
rect 963 752 964 755
rect 774 729 794 733
rect 790 728 794 729
rect 748 717 875 720
rect 881 717 882 720
rect 748 716 882 717
rect 961 704 964 752
rect 727 700 821 703
rect 831 701 974 704
rect 818 696 821 700
rect 770 692 774 693
rect 770 643 774 688
rect 1008 682 1011 962
rect 545 640 774 643
rect 545 639 770 640
rect 1007 630 1011 682
rect 512 626 546 630
rect 601 627 1011 630
rect 1007 626 1011 627
rect 542 622 546 626
rect 542 619 611 622
rect 608 615 611 619
rect 1015 615 1019 970
rect 416 609 504 613
rect 509 609 589 612
rect 608 611 1019 615
rect 1026 601 1029 982
rect 1036 886 1039 995
rect 1170 992 1173 998
rect 1213 998 1239 1001
rect 1243 998 1244 1001
rect 1289 1000 1292 1006
rect 1313 1001 1332 1004
rect 1289 997 1296 1000
rect 1313 996 1316 1001
rect 1336 1002 1375 1003
rect 1336 1000 1371 1002
rect 1163 991 1173 992
rect 1199 991 1218 994
rect 1109 988 1121 991
rect 1163 989 1165 991
rect 1118 924 1121 988
rect 1169 989 1173 991
rect 1181 988 1202 991
rect 1215 988 1263 991
rect 1326 991 1385 994
rect 1296 986 1299 989
rect 1206 971 1209 983
rect 1131 968 1209 971
rect 1296 983 1354 986
rect 1131 939 1134 968
rect 1285 964 1289 982
rect 1166 960 1289 964
rect 1166 934 1170 960
rect 1285 959 1289 960
rect 1300 945 1358 948
rect 1185 940 1267 943
rect 1300 942 1303 945
rect 1330 937 1389 940
rect 1170 930 1191 933
rect 1217 930 1243 933
rect 1247 930 1248 933
rect 1293 931 1300 934
rect 1213 924 1216 930
rect 1118 921 1216 924
rect 1293 925 1296 931
rect 1340 929 1375 931
rect 1340 928 1379 929
rect 1237 922 1296 925
rect 1132 901 1204 903
rect 1128 899 1204 901
rect 1036 883 1151 886
rect 1036 882 1049 883
rect 1200 866 1204 899
rect 1346 892 1349 928
rect 1476 892 1486 893
rect 1346 889 1417 892
rect 1133 863 1213 866
rect 1413 865 1416 889
rect 1476 891 1478 892
rect 1469 887 1478 891
rect 1483 887 1486 892
rect 1469 886 1486 887
rect 1133 857 1136 863
rect 1094 854 1136 857
rect 1209 856 1212 863
rect 1233 861 1292 864
rect 1094 812 1097 854
rect 1166 853 1187 856
rect 1213 853 1239 856
rect 1243 853 1244 856
rect 1289 855 1292 861
rect 1313 856 1332 859
rect 1289 852 1296 855
rect 1313 851 1316 856
rect 1336 857 1375 858
rect 1336 855 1371 857
rect 1109 843 1121 846
rect 1093 746 1097 812
rect 1118 779 1121 843
rect 1181 843 1263 846
rect 1326 846 1385 849
rect 1296 841 1299 844
rect 1296 838 1354 841
rect 1285 819 1289 837
rect 1395 823 1412 826
rect 1474 820 1520 823
rect 1166 815 1289 819
rect 1166 789 1170 815
rect 1285 814 1289 815
rect 1300 800 1358 803
rect 1185 795 1267 798
rect 1300 797 1303 800
rect 1330 792 1389 795
rect 1517 790 1520 820
rect 1532 805 1536 1069
rect 1550 927 1553 1077
rect 1602 1051 1605 1072
rect 1687 1078 1818 1081
rect 1825 1085 1828 1087
rect 1569 1033 1640 1036
rect 1569 945 1572 1033
rect 1637 1029 1640 1033
rect 1565 942 1572 945
rect 1584 980 1623 984
rect 1550 924 1558 927
rect 1555 919 1558 924
rect 1555 916 1565 919
rect 1562 895 1565 916
rect 1557 869 1563 874
rect 1557 864 1558 869
rect 1557 863 1563 864
rect 1532 802 1566 805
rect 1524 790 1553 791
rect 1170 785 1191 788
rect 1217 785 1243 788
rect 1247 785 1248 788
rect 1293 786 1300 789
rect 1213 779 1216 785
rect 1118 776 1216 779
rect 1293 780 1296 786
rect 1340 784 1375 786
rect 1517 787 1553 790
rect 1379 784 1415 786
rect 1340 783 1415 784
rect 1468 786 1472 787
rect 1451 783 1476 786
rect 1237 777 1296 780
rect 1383 755 1387 758
rect 1042 738 1089 741
rect 435 598 1029 601
rect 332 589 355 594
rect 328 587 355 589
rect 224 564 228 584
rect 224 563 595 564
rect 224 562 964 563
rect 224 560 1019 562
rect 224 559 228 560
rect 593 559 1019 560
rect 951 558 1019 559
rect 63 545 413 548
rect 135 526 164 530
rect 71 522 138 526
rect 71 479 76 522
rect 145 515 398 519
rect 35 474 76 479
rect 71 380 76 474
rect 86 457 90 508
rect 145 480 150 515
rect 393 511 397 515
rect 163 502 164 505
rect 168 502 252 505
rect 256 502 345 505
rect 249 484 393 487
rect 144 476 156 480
rect 249 480 252 484
rect 161 476 172 480
rect 301 475 302 478
rect 85 455 90 457
rect 85 419 89 455
rect 229 454 277 457
rect 229 453 286 454
rect 274 450 286 453
rect 299 444 302 475
rect 342 470 345 476
rect 342 467 393 470
rect 408 467 413 545
rect 435 480 438 549
rect 454 491 457 549
rect 466 513 469 549
rect 478 497 479 502
rect 528 501 532 535
rect 570 516 818 520
rect 570 512 574 516
rect 578 504 623 505
rect 627 504 716 507
rect 542 503 545 504
rect 475 478 479 497
rect 540 500 545 503
rect 578 503 716 504
rect 720 503 803 507
rect 578 502 626 503
rect 578 500 581 502
rect 540 497 581 500
rect 475 475 529 478
rect 540 467 545 497
rect 575 486 722 489
rect 719 482 722 486
rect 567 480 574 481
rect 567 478 568 480
rect 561 476 568 478
rect 572 476 574 480
rect 561 475 574 476
rect 623 478 627 481
rect 623 470 626 478
rect 575 467 626 470
rect 719 478 720 482
rect 737 480 756 484
rect 814 482 818 516
rect 1034 494 1037 618
rect 1042 614 1045 738
rect 1086 737 1089 738
rect 1105 738 1148 741
rect 1152 738 1153 741
rect 1105 737 1108 738
rect 1086 734 1108 737
rect 1132 721 1212 724
rect 1132 715 1135 721
rect 1093 712 1135 715
rect 1208 714 1211 721
rect 1232 719 1291 722
rect 1460 720 1463 721
rect 1165 711 1186 714
rect 1199 713 1208 714
rect 1199 709 1202 713
rect 1206 710 1208 713
rect 1212 711 1238 714
rect 1242 711 1243 714
rect 1288 713 1291 719
rect 1312 714 1331 717
rect 1288 710 1295 713
rect 1206 709 1212 710
rect 1312 709 1315 714
rect 1450 717 1463 720
rect 1335 715 1374 716
rect 1335 713 1370 715
rect 1396 711 1415 714
rect 1199 708 1212 709
rect 1108 701 1120 704
rect 1117 637 1120 701
rect 1180 701 1262 704
rect 1325 704 1384 707
rect 1295 699 1298 702
rect 1295 696 1353 699
rect 1284 677 1288 695
rect 1165 673 1288 677
rect 1165 647 1169 673
rect 1284 672 1288 673
rect 1299 658 1357 661
rect 1184 653 1266 656
rect 1299 655 1302 658
rect 1329 650 1388 653
rect 1169 643 1190 646
rect 1216 643 1242 646
rect 1246 643 1247 646
rect 1292 644 1299 647
rect 1212 637 1215 643
rect 1054 633 1106 635
rect 1117 634 1215 637
rect 1292 638 1295 644
rect 1339 642 1374 644
rect 1396 644 1399 711
rect 1378 642 1399 644
rect 1339 641 1399 642
rect 1403 675 1438 679
rect 1236 635 1295 638
rect 1054 632 1102 633
rect 1342 627 1349 628
rect 1342 625 1343 627
rect 1058 622 1343 625
rect 1348 622 1349 627
rect 1342 621 1349 622
rect 1056 617 1063 618
rect 1056 612 1057 617
rect 1062 614 1101 617
rect 1403 617 1406 675
rect 1460 671 1463 717
rect 1412 667 1463 671
rect 1062 612 1063 614
rect 1139 613 1396 616
rect 1400 614 1408 617
rect 1056 611 1063 612
rect 1412 606 1417 667
rect 1072 604 1077 605
rect 1071 603 1113 604
rect 1412 603 1415 606
rect 1427 603 1458 607
rect 1071 600 1415 603
rect 1071 597 1076 600
rect 1072 595 1076 597
rect 1042 573 1062 577
rect 1042 564 1046 573
rect 1064 558 1066 564
rect 1061 517 1066 558
rect 800 478 808 482
rect 813 480 818 482
rect 813 478 1040 480
rect 408 462 545 467
rect 410 461 419 462
rect 620 459 623 467
rect 547 456 558 458
rect 620 456 634 459
rect 547 455 552 456
rect 328 452 552 455
rect 556 452 558 456
rect 328 451 558 452
rect 658 450 661 477
rect 720 468 723 478
rect 814 477 1040 478
rect 827 476 1040 477
rect 1026 468 1030 469
rect 720 464 1030 468
rect 673 456 732 459
rect 563 447 661 450
rect 760 456 1022 459
rect 746 452 750 455
rect 746 449 813 452
rect 251 443 304 444
rect 169 440 304 443
rect 563 442 567 447
rect 169 434 172 440
rect 118 431 183 434
rect 85 415 126 419
rect 122 408 126 415
rect 75 376 76 380
rect 83 406 86 407
rect 83 403 90 406
rect 83 338 86 403
rect 126 404 159 407
rect 179 407 182 431
rect 261 431 346 434
rect 350 431 371 434
rect 447 433 512 436
rect 315 426 364 427
rect 315 424 360 426
rect 315 415 318 424
rect 230 403 263 406
rect 243 399 246 403
rect 355 399 358 405
rect 243 396 358 399
rect 319 387 320 390
rect 317 339 320 387
rect 368 381 371 431
rect 508 430 512 433
rect 563 430 566 442
rect 809 439 813 449
rect 570 436 590 438
rect 570 435 586 436
rect 570 431 571 435
rect 575 432 586 435
rect 590 433 675 436
rect 774 436 839 439
rect 575 431 590 432
rect 570 430 578 431
rect 508 427 566 430
rect 412 405 419 408
rect 362 377 396 381
rect 356 376 396 377
rect 83 335 177 338
rect 187 336 330 339
rect 174 331 177 335
rect 346 331 350 363
rect 349 328 350 331
rect 325 305 356 309
rect 306 304 330 305
rect 263 301 330 304
rect 263 300 266 301
rect 207 297 266 300
rect 207 288 211 297
rect 117 285 211 288
rect 82 257 89 260
rect 82 192 85 257
rect 125 258 158 261
rect 178 261 181 285
rect 260 285 345 288
rect 314 279 317 281
rect 314 276 361 279
rect 139 223 142 258
rect 229 257 262 260
rect 242 253 245 257
rect 354 253 357 259
rect 242 250 357 253
rect 318 241 319 244
rect 239 225 242 241
rect 139 219 232 223
rect 238 222 305 225
rect 227 206 232 219
rect 227 202 300 206
rect 316 193 319 241
rect 369 237 372 376
rect 380 353 401 357
rect 412 340 415 405
rect 455 406 488 409
rect 508 409 511 427
rect 647 425 805 428
rect 731 418 790 421
rect 473 357 477 406
rect 559 405 592 408
rect 572 401 575 405
rect 684 401 687 407
rect 572 398 687 401
rect 731 399 735 418
rect 703 395 735 399
rect 739 408 746 411
rect 648 389 649 392
rect 486 365 487 368
rect 492 365 583 368
rect 646 341 649 389
rect 689 379 723 383
rect 683 378 723 379
rect 672 361 676 365
rect 412 337 506 340
rect 516 338 649 341
rect 673 337 676 361
rect 699 350 727 353
rect 739 343 742 408
rect 782 409 815 412
rect 835 412 838 436
rect 917 436 1002 439
rect 894 428 968 430
rect 894 427 972 428
rect 788 362 791 393
rect 760 359 791 362
rect 798 354 802 409
rect 886 408 919 411
rect 899 404 902 408
rect 1011 404 1014 410
rect 899 401 1014 404
rect 807 367 810 392
rect 975 392 976 395
rect 824 355 883 358
rect 891 354 895 392
rect 973 344 976 392
rect 739 340 833 343
rect 843 341 986 344
rect 503 333 506 337
rect 830 336 833 340
rect 380 325 486 329
rect 781 329 785 330
rect 720 327 785 329
rect 801 329 821 332
rect 801 327 804 329
rect 561 326 804 327
rect 561 324 724 326
rect 781 324 804 326
rect 818 328 821 329
rect 881 329 929 332
rect 818 324 820 328
rect 824 324 825 327
rect 561 308 564 324
rect 729 318 730 322
rect 734 318 739 321
rect 729 317 739 318
rect 743 317 748 321
rect 881 320 884 329
rect 812 318 884 320
rect 808 317 884 318
rect 890 311 895 314
rect 381 305 564 308
rect 590 307 895 311
rect 590 306 713 307
rect 591 290 596 306
rect 923 293 926 329
rect 1007 312 1015 315
rect 446 287 511 290
rect 380 276 404 279
rect 400 256 404 276
rect 478 271 481 287
rect 411 259 418 262
rect 400 253 406 256
rect 364 236 394 237
rect 364 231 393 236
rect 334 202 354 206
rect 82 189 176 192
rect 186 190 329 193
rect 173 185 176 189
rect 340 178 355 181
rect 365 116 371 231
rect 403 215 406 253
rect 392 206 396 207
rect 380 202 396 206
rect 376 169 380 178
rect 392 181 396 202
rect 411 194 414 259
rect 454 260 487 263
rect 507 263 510 287
rect 589 287 674 290
rect 773 290 838 293
rect 716 282 794 285
rect 717 273 721 282
rect 798 282 800 285
rect 647 270 721 273
rect 427 207 431 223
rect 454 217 464 219
rect 454 215 459 217
rect 458 211 459 215
rect 458 210 464 211
rect 469 213 472 260
rect 558 259 591 262
rect 571 255 574 259
rect 683 255 686 261
rect 571 252 686 255
rect 738 262 745 265
rect 478 247 481 248
rect 647 243 648 246
rect 478 221 481 243
rect 493 225 631 228
rect 469 209 568 213
rect 645 195 648 243
rect 687 233 723 236
rect 661 209 720 214
rect 738 197 741 262
rect 781 263 814 266
rect 834 266 837 290
rect 916 290 1001 293
rect 1011 284 1015 312
rect 971 281 1015 284
rect 971 277 974 281
rect 792 236 796 250
rect 765 232 796 236
rect 765 222 769 232
rect 792 231 796 232
rect 801 227 805 263
rect 885 262 918 265
rect 898 258 901 262
rect 1010 258 1013 264
rect 898 255 1013 258
rect 974 246 975 249
rect 785 223 805 227
rect 801 222 805 223
rect 746 218 769 222
rect 746 205 750 218
rect 759 211 886 214
rect 892 211 893 214
rect 759 210 893 211
rect 746 201 797 205
rect 972 198 975 246
rect 993 224 1001 226
rect 993 220 995 224
rect 1000 220 1001 224
rect 993 218 1001 220
rect 411 191 505 194
rect 515 192 658 195
rect 712 194 725 196
rect 738 194 832 197
rect 842 195 985 198
rect 950 194 963 195
rect 502 187 505 191
rect 680 193 725 194
rect 680 192 724 193
rect 680 190 717 192
rect 721 188 724 192
rect 829 190 832 194
rect 721 186 770 188
rect 721 184 762 186
rect 392 177 469 181
rect 466 173 469 177
rect 549 176 551 181
rect 760 180 762 184
rect 767 184 770 186
rect 781 186 785 187
rect 767 180 769 184
rect 729 176 730 179
rect 760 178 769 180
rect 797 182 800 184
rect 549 173 554 176
rect 376 168 428 169
rect 376 165 432 168
rect 450 144 454 169
rect 466 169 554 173
rect 466 168 469 169
rect 729 158 734 176
rect 729 155 766 158
rect 731 154 766 155
rect 647 153 652 154
rect 781 137 785 182
rect 556 134 785 137
rect 556 133 781 134
rect 797 132 800 177
rect 950 170 952 176
rect 958 170 959 176
rect 950 168 959 170
rect 879 133 886 137
rect 993 133 997 218
rect 1019 176 1022 456
rect 879 132 997 133
rect 797 129 997 132
rect 1018 124 1022 176
rect 523 120 557 124
rect 612 121 1022 124
rect 1018 120 1022 121
rect 553 116 557 120
rect 365 88 368 116
rect 553 113 622 116
rect 619 109 622 113
rect 1026 109 1030 464
rect 379 104 422 107
rect 427 103 515 107
rect 520 103 600 106
rect 619 105 1030 109
rect 1037 95 1040 476
rect 1062 443 1066 517
rect 1072 411 1077 595
rect 1174 594 1178 595
rect 1096 593 1305 594
rect 1468 593 1472 783
rect 1096 590 1472 593
rect 1152 573 1155 583
rect 1096 548 1100 566
rect 1096 546 1142 548
rect 1096 545 1146 546
rect 1152 517 1155 568
rect 1174 564 1178 590
rect 1227 589 1472 590
rect 1355 588 1472 589
rect 1532 773 1554 777
rect 1343 567 1344 571
rect 1348 567 1508 571
rect 1228 561 1237 562
rect 1228 558 1471 561
rect 1174 556 1178 557
rect 1154 497 1234 500
rect 1154 491 1157 497
rect 1230 492 1233 497
rect 1254 495 1313 498
rect 446 92 1040 95
rect 1045 406 1077 411
rect 1045 193 1048 406
rect 1062 375 1066 392
rect 1083 390 1087 489
rect 1115 488 1157 491
rect 1224 490 1235 492
rect 1187 487 1208 490
rect 1224 486 1225 490
rect 1229 486 1230 490
rect 1234 487 1260 490
rect 1234 486 1235 487
rect 1264 487 1265 490
rect 1310 489 1313 495
rect 1334 490 1353 493
rect 1310 486 1317 489
rect 1224 484 1235 486
rect 1334 485 1337 490
rect 1357 491 1396 492
rect 1357 489 1392 491
rect 1130 477 1142 480
rect 1139 413 1142 477
rect 1202 477 1284 480
rect 1347 480 1406 483
rect 1317 475 1320 478
rect 1317 472 1375 475
rect 1466 473 1469 558
rect 1306 453 1310 471
rect 1466 468 1489 473
rect 1187 449 1310 453
rect 1187 423 1191 449
rect 1306 448 1310 449
rect 1455 438 1490 441
rect 1455 437 1495 438
rect 1321 434 1379 437
rect 1206 429 1288 432
rect 1321 431 1324 434
rect 1351 426 1410 429
rect 1191 419 1212 422
rect 1238 419 1264 422
rect 1268 419 1269 422
rect 1314 420 1321 423
rect 1234 413 1237 419
rect 1139 410 1237 413
rect 1314 414 1317 420
rect 1361 418 1396 420
rect 1503 420 1508 567
rect 1532 443 1536 773
rect 1563 755 1566 802
rect 1570 802 1573 932
rect 1584 818 1588 980
rect 1638 967 1641 993
rect 1665 983 1668 1001
rect 1596 964 1641 967
rect 1596 828 1599 964
rect 1638 960 1641 964
rect 1603 814 1606 951
rect 1665 940 1668 979
rect 1687 976 1690 1078
rect 1825 1070 1829 1085
rect 1720 1067 1829 1070
rect 1687 973 1695 976
rect 1692 948 1695 973
rect 1641 937 1668 940
rect 1665 936 1668 937
rect 1675 945 1695 948
rect 1704 961 1707 1046
rect 1720 1017 1723 1067
rect 1733 1055 1742 1058
rect 1704 948 1707 957
rect 1704 945 1723 948
rect 1675 929 1678 945
rect 1652 926 1678 929
rect 1682 938 1703 941
rect 1637 876 1640 889
rect 1652 877 1655 926
rect 1682 882 1685 938
rect 1720 933 1723 945
rect 1708 930 1723 933
rect 1732 946 1735 963
rect 1739 946 1742 1055
rect 1799 1020 1802 1030
rect 1748 1019 1802 1020
rect 1751 1017 1802 1019
rect 1732 943 1742 946
rect 1732 930 1735 943
rect 1750 938 1768 941
rect 1708 898 1711 930
rect 1630 873 1640 876
rect 1570 800 1621 802
rect 1570 799 1624 800
rect 1603 779 1606 788
rect 1573 776 1606 779
rect 1561 752 1569 755
rect 1553 670 1557 727
rect 1566 716 1569 752
rect 1573 685 1576 776
rect 1630 764 1633 873
rect 1637 856 1640 873
rect 1647 874 1655 877
rect 1665 879 1685 882
rect 1696 895 1711 898
rect 1647 804 1650 874
rect 1665 862 1668 879
rect 1665 773 1668 858
rect 1696 772 1699 895
rect 1799 887 1802 1017
rect 1808 994 1819 997
rect 1808 989 1812 994
rect 1817 989 1819 994
rect 1808 986 1819 989
rect 1812 982 1819 986
rect 1808 979 1819 982
rect 1825 965 1829 1067
rect 1819 960 1829 965
rect 1819 953 1820 960
rect 1825 953 1829 960
rect 1819 950 1829 953
rect 1704 882 1707 883
rect 1704 879 1731 882
rect 1704 839 1707 879
rect 1800 874 1807 877
rect 1731 841 1734 859
rect 1704 835 1715 839
rect 1704 818 1707 835
rect 1712 785 1715 835
rect 1731 838 1787 841
rect 1731 826 1734 838
rect 1732 786 1735 790
rect 1800 786 1803 874
rect 1838 871 1841 1087
rect 1883 1067 1887 1115
rect 1916 1105 1917 1111
rect 1873 1062 1887 1067
rect 1838 869 1853 871
rect 1838 861 1844 869
rect 1850 861 1853 869
rect 1838 860 1853 861
rect 1808 858 1853 860
rect 1808 857 1841 858
rect 1808 813 1811 857
rect 1807 810 1812 813
rect 1712 782 1721 785
rect 1732 783 1803 786
rect 1696 768 1713 772
rect 1630 761 1639 764
rect 1709 749 1713 768
rect 1581 744 1713 749
rect 1581 689 1584 744
rect 1718 717 1721 782
rect 1733 775 1769 776
rect 1733 771 1760 775
rect 1733 728 1741 771
rect 1768 771 1769 775
rect 1809 745 1812 810
rect 1772 742 1812 745
rect 1817 736 1820 836
rect 1816 731 1869 736
rect 1740 722 1741 728
rect 1595 712 1678 716
rect 1718 714 1781 717
rect 1568 682 1576 685
rect 1549 666 1557 670
rect 1571 673 1642 676
rect 1532 433 1536 437
rect 1549 434 1552 666
rect 1571 585 1574 673
rect 1639 669 1642 673
rect 1567 582 1574 585
rect 1400 418 1437 420
rect 1361 417 1437 418
rect 1258 411 1317 414
rect 1083 389 1276 390
rect 1083 388 1332 389
rect 1083 385 1419 388
rect 1062 372 1171 375
rect 1062 371 1066 372
rect 1152 352 1232 355
rect 1152 346 1155 352
rect 1113 343 1155 346
rect 1228 345 1231 352
rect 1252 350 1311 353
rect 1185 342 1206 345
rect 1222 341 1223 345
rect 1227 341 1228 345
rect 1232 342 1258 345
rect 1262 342 1263 345
rect 1308 344 1311 350
rect 1332 345 1351 348
rect 1308 341 1315 344
rect 1222 339 1231 341
rect 1332 340 1335 345
rect 1355 346 1394 347
rect 1355 344 1390 346
rect 1128 332 1140 335
rect 1137 268 1140 332
rect 1200 332 1282 335
rect 1345 335 1404 338
rect 1315 330 1318 333
rect 1315 327 1373 330
rect 1304 308 1308 326
rect 1416 316 1419 385
rect 1185 304 1308 308
rect 1185 278 1189 304
rect 1304 303 1308 304
rect 1365 313 1419 316
rect 1433 317 1437 417
rect 1503 416 1515 420
rect 1511 332 1515 416
rect 1548 369 1552 434
rect 1572 442 1575 572
rect 1581 544 1584 659
rect 1622 649 1635 652
rect 1622 647 1625 649
rect 1599 644 1625 647
rect 1589 623 1623 627
rect 1589 461 1593 623
rect 1632 616 1635 649
rect 1631 612 1635 616
rect 1640 607 1643 633
rect 1667 627 1670 641
rect 1654 623 1670 627
rect 1600 603 1643 607
rect 1600 454 1604 603
rect 1640 600 1643 603
rect 1614 592 1617 595
rect 1649 592 1652 608
rect 1614 589 1652 592
rect 1614 521 1617 589
rect 1667 580 1670 623
rect 1643 577 1670 580
rect 1667 576 1670 577
rect 1675 568 1678 712
rect 1778 711 1781 714
rect 1778 708 1856 711
rect 1722 705 1770 706
rect 1722 703 1767 705
rect 1706 601 1709 686
rect 1722 659 1725 703
rect 1735 695 1744 698
rect 1706 588 1709 597
rect 1706 585 1725 588
rect 1656 565 1678 568
rect 1684 578 1705 581
rect 1614 520 1627 521
rect 1614 517 1624 520
rect 1639 516 1642 529
rect 1632 513 1642 516
rect 1572 440 1623 442
rect 1572 439 1626 440
rect 1572 429 1575 439
rect 1632 404 1635 513
rect 1639 496 1642 513
rect 1649 444 1652 516
rect 1656 506 1659 565
rect 1684 522 1687 578
rect 1722 573 1725 585
rect 1710 570 1725 573
rect 1734 586 1737 603
rect 1741 586 1744 695
rect 1801 660 1804 670
rect 1750 659 1804 660
rect 1753 657 1804 659
rect 1734 583 1744 586
rect 1734 570 1737 583
rect 1752 578 1770 581
rect 1710 538 1713 570
rect 1667 519 1687 522
rect 1698 535 1713 538
rect 1656 502 1660 506
rect 1667 502 1670 519
rect 1632 401 1641 404
rect 1657 388 1660 502
rect 1667 413 1670 498
rect 1698 412 1701 535
rect 1801 527 1804 657
rect 1706 522 1709 523
rect 1706 519 1733 522
rect 1706 486 1709 519
rect 1802 514 1809 517
rect 1784 502 1796 506
rect 1706 483 1723 486
rect 1706 458 1709 483
rect 1698 408 1715 412
rect 1657 385 1666 388
rect 1542 367 1552 369
rect 1542 361 1544 367
rect 1550 363 1552 367
rect 1550 361 1551 363
rect 1542 360 1551 361
rect 1565 348 1646 353
rect 1514 328 1515 332
rect 1599 325 1603 334
rect 1599 324 1600 325
rect 1517 320 1600 324
rect 1639 323 1646 348
rect 1663 347 1666 385
rect 1685 355 1690 398
rect 1711 391 1715 408
rect 1720 357 1723 483
rect 1733 483 1736 499
rect 1778 495 1786 502
rect 1791 495 1796 502
rect 1778 493 1796 495
rect 1733 480 1782 483
rect 1733 466 1736 480
rect 1734 426 1737 430
rect 1802 426 1805 514
rect 1824 478 1844 482
rect 1820 477 1844 478
rect 1734 423 1805 426
rect 1735 415 1771 416
rect 1735 411 1762 415
rect 1735 368 1743 411
rect 1770 411 1771 415
rect 1765 384 1796 388
rect 1810 387 1814 431
rect 1742 362 1743 368
rect 1720 354 1772 357
rect 1663 346 1681 347
rect 1709 346 1766 349
rect 1663 342 1713 346
rect 1663 323 1667 324
rect 1433 314 1444 317
rect 1448 314 1453 317
rect 1489 315 1493 316
rect 1365 302 1368 313
rect 1415 306 1432 309
rect 1429 298 1432 306
rect 1429 294 1435 298
rect 1489 297 1493 309
rect 1439 294 1440 297
rect 1489 294 1506 297
rect 1319 289 1377 292
rect 1204 284 1286 287
rect 1319 286 1322 289
rect 1517 287 1521 320
rect 1599 319 1603 320
rect 1639 316 1667 323
rect 1349 281 1408 284
rect 1511 283 1520 287
rect 1189 274 1210 277
rect 1236 274 1262 277
rect 1266 274 1267 277
rect 1312 275 1319 278
rect 1232 268 1235 274
rect 1137 265 1235 268
rect 1312 269 1315 275
rect 1359 273 1394 275
rect 1398 273 1436 275
rect 1359 272 1436 273
rect 1256 266 1315 269
rect 1355 253 1419 256
rect 1084 252 1099 253
rect 1089 251 1099 252
rect 1089 250 1306 251
rect 1355 250 1358 253
rect 1089 248 1358 250
rect 1084 247 1358 248
rect 1063 232 1067 233
rect 1063 229 1170 232
rect 1063 193 1067 229
rect 1365 218 1368 245
rect 1153 210 1233 213
rect 1153 204 1156 210
rect 1229 205 1232 210
rect 1253 208 1312 211
rect 1114 201 1156 204
rect 1222 204 1232 205
rect 1168 199 1182 202
rect 1186 200 1207 203
rect 1186 199 1188 200
rect 1222 200 1223 204
rect 1227 203 1232 204
rect 1227 200 1229 203
rect 1222 199 1229 200
rect 1233 200 1259 203
rect 1263 200 1264 203
rect 1309 202 1312 208
rect 1333 203 1352 206
rect 1309 199 1316 202
rect 1045 190 1069 193
rect 1129 190 1141 193
rect 1045 131 1048 190
rect 1114 153 1116 157
rect 1045 128 1052 131
rect 1111 131 1115 153
rect 1056 128 1115 131
rect 1045 91 1048 128
rect 1138 126 1141 190
rect 1168 188 1171 199
rect 1333 198 1336 203
rect 1356 204 1395 205
rect 1356 202 1391 204
rect 1201 190 1283 193
rect 1346 193 1405 196
rect 1316 188 1319 191
rect 1149 185 1171 188
rect 1149 158 1152 185
rect 1316 185 1374 188
rect 1305 166 1309 184
rect 1416 181 1419 253
rect 1433 227 1436 272
rect 1433 224 1447 227
rect 1451 224 1456 227
rect 1492 221 1504 224
rect 1512 181 1515 283
rect 1365 175 1366 179
rect 1416 178 1516 181
rect 1416 175 1419 178
rect 1186 162 1309 166
rect 1186 136 1190 162
rect 1305 161 1309 162
rect 1363 162 1366 175
rect 1544 174 1549 301
rect 1639 288 1645 294
rect 1639 285 1650 288
rect 1639 284 1649 285
rect 1639 278 1640 284
rect 1646 278 1649 284
rect 1639 276 1649 278
rect 1646 226 1659 228
rect 1646 224 1652 226
rect 1646 220 1647 224
rect 1651 220 1652 224
rect 1657 220 1659 226
rect 1646 217 1659 220
rect 1451 166 1454 173
rect 1416 163 1454 166
rect 1363 160 1368 162
rect 1363 158 1364 160
rect 1320 147 1378 150
rect 1205 142 1287 145
rect 1320 144 1323 147
rect 1350 139 1409 142
rect 1434 139 1440 142
rect 1444 139 1457 142
rect 1190 132 1211 135
rect 1237 132 1263 135
rect 1267 132 1268 135
rect 1313 133 1320 136
rect 1233 126 1236 132
rect 1138 123 1236 126
rect 1313 127 1316 133
rect 1360 131 1395 133
rect 1360 130 1399 131
rect 1257 124 1316 127
rect 1388 126 1391 130
rect 1434 126 1437 139
rect 1492 135 1534 139
rect 1388 123 1437 126
rect 1497 112 1502 113
rect 1497 106 1498 112
rect 1364 101 1365 105
rect 1098 95 1102 96
rect 365 81 366 88
rect 668 83 669 87
rect 673 85 676 87
rect 673 83 1047 85
rect 668 82 1047 83
rect 950 46 954 52
rect 959 46 983 52
rect 950 44 983 46
rect 1039 36 1042 82
rect 1098 61 1102 90
rect 1097 60 1238 61
rect 1097 56 1349 60
rect 1038 29 1056 36
rect 1039 27 1042 29
rect 1364 22 1367 101
rect 1364 18 1398 22
rect 1403 18 1410 22
rect 1497 8 1503 106
rect 1544 48 1547 174
rect 1580 91 1581 97
rect 1580 53 1584 91
rect 1630 86 1636 88
rect 1633 79 1636 86
rect 1534 43 1547 48
rect 1578 51 1588 53
rect 1578 44 1581 51
rect 1586 44 1588 51
rect 1630 49 1636 79
rect 1650 62 1654 77
rect 1578 42 1588 44
rect 1625 45 1637 49
rect 1625 39 1627 45
rect 1633 39 1637 45
rect 1625 37 1637 39
rect 1663 33 1667 316
rect 1698 245 1701 330
rect 1709 303 1713 342
rect 1727 339 1736 342
rect 1709 300 1710 303
rect 1726 230 1729 247
rect 1733 230 1736 339
rect 1763 311 1766 346
rect 1793 322 1796 384
rect 1826 357 1830 358
rect 1805 354 1830 357
rect 1777 318 1796 322
rect 1763 308 1818 311
rect 1742 303 1796 304
rect 1745 301 1796 303
rect 1780 281 1783 289
rect 1769 278 1783 281
rect 1769 250 1772 278
rect 1726 227 1736 230
rect 1726 214 1729 227
rect 1745 220 1772 224
rect 1698 166 1701 167
rect 1698 163 1725 166
rect 1698 102 1701 163
rect 1743 155 1747 220
rect 1754 213 1757 216
rect 1754 210 1761 213
rect 1754 162 1757 210
rect 1769 206 1772 220
rect 1768 203 1772 206
rect 1768 167 1771 203
rect 1793 178 1796 301
rect 1790 175 1796 178
rect 1790 174 1793 175
rect 1776 171 1793 174
rect 1801 167 1819 171
rect 1754 159 1764 162
rect 1779 160 1786 163
rect 1743 152 1775 155
rect 1743 151 1771 152
rect 1725 127 1728 143
rect 1705 124 1728 127
rect 1678 77 1679 81
rect 1676 56 1679 77
rect 1676 52 1696 56
rect 1663 30 1697 33
rect 1625 26 1645 30
rect 1523 18 1683 22
rect 1706 12 1709 124
rect 1725 110 1728 124
rect 1744 92 1747 135
rect 1718 89 1747 92
rect 1718 34 1721 89
rect 1768 87 1771 151
rect 1779 116 1782 160
rect 1816 158 1819 167
rect 1794 155 1819 158
rect 1779 112 1783 116
rect 1726 70 1729 74
rect 1794 70 1797 155
rect 1726 67 1797 70
rect 1736 37 1740 52
rect 1786 53 1795 55
rect 1786 49 1787 53
rect 1791 50 1795 53
rect 1799 50 1800 55
rect 1791 49 1799 50
rect 1786 48 1799 49
rect 1809 34 1812 141
rect 1718 14 1721 29
rect 1759 27 1761 31
rect 1765 27 1772 31
rect 1759 26 1772 27
rect 1802 31 1812 34
rect 1759 24 1775 26
rect 1809 20 1812 31
rect 1496 7 1517 8
rect 1496 5 1660 7
rect 1826 5 1830 354
rect 1838 22 1844 477
rect 1851 271 1856 708
rect 1863 548 1869 731
rect 1863 482 1870 548
rect 1843 18 1844 22
rect 1850 10 1856 271
rect 1864 21 1870 482
rect 1874 280 1878 1062
rect 1894 995 1903 998
rect 1894 991 1895 995
rect 1899 991 1903 995
rect 1894 989 1903 991
rect 1908 989 1909 998
rect 1884 963 1893 965
rect 1884 961 1898 963
rect 1884 955 1886 961
rect 1894 955 1898 961
rect 1914 959 1917 1105
rect 1925 1097 1944 1100
rect 1926 1082 2006 1086
rect 1952 975 2708 978
rect 2712 975 2803 978
rect 2800 970 2803 975
rect 1933 965 1956 966
rect 1933 963 2708 965
rect 1953 962 2708 963
rect 1884 946 1898 955
rect 1912 958 1930 959
rect 1912 955 2882 958
rect 1912 954 1964 955
rect 1914 953 1917 954
rect 1889 944 1898 946
rect 1951 947 1956 948
rect 1951 944 2655 947
rect 1893 599 1897 944
rect 1906 914 1912 915
rect 1951 914 1956 944
rect 1906 912 1956 914
rect 1906 910 1955 912
rect 1906 776 1912 910
rect 2005 854 2009 924
rect 2084 894 2088 895
rect 2087 889 2088 894
rect 2084 823 2088 889
rect 2211 852 2214 888
rect 2288 827 2292 924
rect 2493 905 2496 909
rect 2340 901 2483 904
rect 2493 902 2587 905
rect 2350 882 2353 901
rect 2455 892 2570 895
rect 2349 879 2353 882
rect 2384 879 2510 882
rect 2350 853 2353 879
rect 2384 869 2429 872
rect 2426 855 2429 869
rect 2350 850 2351 853
rect 2426 852 2490 855
rect 2312 841 2427 844
rect 2312 835 2315 841
rect 2424 837 2427 841
rect 2487 837 2490 852
rect 2407 834 2440 837
rect 2288 824 2354 827
rect 1932 822 1945 823
rect 1932 813 1934 822
rect 1942 813 1945 822
rect 2084 820 2131 823
rect 1932 806 1945 813
rect 2324 806 2409 809
rect 2488 809 2491 833
rect 2507 836 2510 879
rect 2511 833 2544 836
rect 2584 837 2587 902
rect 2632 903 2635 935
rect 2652 922 2655 944
rect 2652 919 2788 922
rect 2800 914 2803 945
rect 2878 928 2881 955
rect 2800 911 2807 914
rect 2853 907 2856 911
rect 2711 903 2843 906
rect 2853 904 2947 907
rect 2632 900 2674 903
rect 2600 892 2660 895
rect 2580 834 2587 837
rect 2413 806 2433 809
rect 2487 806 2552 809
rect 1932 803 2257 806
rect 1932 802 2128 803
rect 2140 802 2203 803
rect 1932 801 2119 802
rect 2141 801 2203 802
rect 2219 801 2257 803
rect 1932 800 1945 801
rect 2123 796 2132 798
rect 1962 795 2132 796
rect 1962 794 2136 795
rect 1962 792 2126 794
rect 2211 793 2215 795
rect 1963 781 1966 792
rect 2211 786 2214 793
rect 1911 771 1912 776
rect 2013 775 2078 778
rect 1944 767 2055 770
rect 2074 759 2077 775
rect 2156 775 2241 778
rect 2254 766 2257 801
rect 2430 792 2433 806
rect 2266 786 2309 791
rect 2430 789 2492 792
rect 2319 775 2449 778
rect 2254 762 2265 766
rect 1909 756 2077 759
rect 1909 639 1912 756
rect 1978 747 1985 750
rect 1908 633 1912 639
rect 1961 632 1965 743
rect 1978 682 1981 747
rect 2021 748 2054 751
rect 2074 751 2077 756
rect 2125 747 2158 750
rect 2138 743 2141 747
rect 2250 743 2253 749
rect 2261 751 2265 762
rect 2319 765 2323 775
rect 2369 767 2434 770
rect 2302 761 2323 765
rect 2261 748 2390 751
rect 2430 753 2433 767
rect 2446 766 2449 775
rect 2489 771 2492 789
rect 2496 767 2508 770
rect 2446 763 2484 766
rect 2406 750 2433 753
rect 2481 754 2484 763
rect 2496 754 2499 767
rect 2512 767 2597 770
rect 2655 767 2660 892
rect 2711 855 2714 903
rect 2722 895 2807 898
rect 2767 887 2868 890
rect 2780 878 2850 881
rect 2780 855 2783 878
rect 2788 865 2791 870
rect 2788 862 2851 865
rect 2672 843 2787 846
rect 2672 837 2675 843
rect 2784 839 2787 843
rect 2848 839 2851 862
rect 2767 836 2800 839
rect 2878 838 2881 894
rect 2716 824 2787 827
rect 2684 808 2769 811
rect 2848 811 2851 835
rect 2871 835 2904 838
rect 2878 834 2881 835
rect 2944 839 2947 904
rect 2955 887 2985 890
rect 2955 878 2985 881
rect 2940 836 2947 839
rect 2773 808 2793 811
rect 2847 808 2912 811
rect 2790 794 2793 808
rect 2790 791 2852 794
rect 2679 777 2809 780
rect 2679 767 2683 777
rect 2729 769 2794 772
rect 2655 763 2683 767
rect 2481 751 2499 754
rect 2751 756 2754 769
rect 2138 740 2253 743
rect 2279 734 2327 741
rect 2214 731 2215 734
rect 2273 733 2327 734
rect 2131 708 2135 731
rect 1998 705 2135 708
rect 2212 683 2215 731
rect 2322 714 2327 733
rect 1978 679 2072 682
rect 2082 680 2215 683
rect 2295 683 2299 711
rect 2326 706 2327 714
rect 2322 705 2327 706
rect 2334 739 2341 742
rect 2230 680 2299 683
rect 2069 675 2072 679
rect 2334 674 2337 739
rect 2387 743 2390 748
rect 2377 740 2410 743
rect 2430 743 2433 750
rect 2570 749 2623 752
rect 2481 739 2514 742
rect 2494 735 2497 739
rect 2606 735 2609 741
rect 2494 732 2609 735
rect 2402 690 2405 732
rect 2489 706 2492 724
rect 2570 723 2571 726
rect 2568 675 2571 723
rect 2334 671 2428 674
rect 2438 672 2581 675
rect 2019 640 2023 644
rect 2023 636 2027 640
rect 2065 638 2068 663
rect 2425 667 2428 671
rect 2298 662 2342 666
rect 2261 643 2268 644
rect 2261 639 2262 643
rect 2266 641 2268 643
rect 2266 639 2272 641
rect 2261 638 2272 639
rect 1961 629 1994 632
rect 2403 624 2406 658
rect 2620 629 2623 749
rect 2639 736 2687 743
rect 2633 735 2687 736
rect 2682 716 2687 735
rect 2686 708 2687 716
rect 2682 707 2687 708
rect 2694 741 2701 744
rect 2694 676 2697 741
rect 2737 742 2770 745
rect 2790 745 2793 769
rect 2806 768 2809 777
rect 2849 773 2852 791
rect 2856 769 2868 772
rect 2806 765 2844 768
rect 2841 756 2844 765
rect 2856 756 2859 769
rect 2872 769 2957 772
rect 2841 753 2859 756
rect 2929 751 2989 754
rect 2763 735 2766 742
rect 2841 741 2874 744
rect 2854 737 2857 741
rect 2966 737 2969 743
rect 2854 734 2969 737
rect 2752 700 2755 731
rect 2763 686 2766 731
rect 2849 708 2852 726
rect 2930 725 2931 728
rect 2928 677 2931 725
rect 2694 673 2788 676
rect 2798 674 2941 677
rect 2785 669 2788 673
rect 2753 662 2754 663
rect 2753 635 2757 662
rect 1917 619 1927 624
rect 1935 619 2406 624
rect 2753 610 2758 635
rect 1920 606 2758 610
rect 2764 599 2767 661
rect 1893 596 2767 599
rect 1893 595 1932 596
rect 2022 589 2028 591
rect 2022 585 2023 589
rect 2027 588 2028 589
rect 2027 585 2034 588
rect 2022 584 2028 585
rect 2261 581 2267 583
rect 2261 577 2262 581
rect 2266 577 2267 581
rect 2224 572 2231 573
rect 1934 568 2231 572
rect 1952 544 2050 546
rect 1952 542 2188 544
rect 1952 538 2182 542
rect 2186 538 2188 542
rect 2042 537 2188 538
rect 2010 521 2110 522
rect 1908 517 2104 521
rect 2108 517 2110 521
rect 1908 516 2110 517
rect 2224 512 2231 568
rect 2261 571 2267 577
rect 2261 567 2262 571
rect 2266 567 2267 571
rect 2261 566 2267 567
rect 2224 511 2916 512
rect 2224 507 2909 511
rect 2913 507 2916 511
rect 2224 506 2916 507
rect 2251 490 2296 493
rect 1981 481 1985 484
rect 1981 476 1982 481
rect 1981 462 1985 476
rect 2197 461 2202 477
rect 2000 455 2029 459
rect 1936 454 1975 455
rect 1994 454 2003 455
rect 1936 451 2003 454
rect 1901 442 1912 443
rect 1901 435 1904 442
rect 1909 437 1912 442
rect 1936 437 1941 451
rect 2010 444 2263 448
rect 1909 435 1941 437
rect 1901 432 1941 435
rect 1913 422 1915 428
rect 1897 224 1901 414
rect 1913 394 1919 422
rect 1913 388 1918 394
rect 1912 264 1918 388
rect 1936 309 1941 432
rect 1951 386 1955 437
rect 1995 418 1999 432
rect 1967 413 2000 418
rect 1995 412 1999 413
rect 2010 409 2015 444
rect 2258 440 2262 444
rect 2028 431 2029 434
rect 2033 431 2117 434
rect 2121 431 2210 434
rect 2293 432 2296 490
rect 2393 430 2397 464
rect 2435 445 2683 449
rect 2435 441 2439 445
rect 2492 433 2581 436
rect 2490 432 2581 433
rect 2585 432 2606 436
rect 2610 432 2668 436
rect 2114 413 2258 416
rect 2440 415 2587 418
rect 2009 405 2021 409
rect 2114 409 2117 413
rect 2584 411 2587 415
rect 2026 405 2037 409
rect 2166 404 2167 407
rect 1950 384 1955 386
rect 1950 348 1954 384
rect 2094 383 2142 386
rect 2094 382 2151 383
rect 2139 379 2151 382
rect 2164 373 2167 404
rect 2178 405 2188 408
rect 2178 400 2180 405
rect 2184 400 2188 405
rect 2178 398 2188 400
rect 2207 399 2210 405
rect 2488 407 2492 410
rect 2179 376 2183 398
rect 2207 396 2258 399
rect 2488 399 2491 407
rect 2440 396 2491 399
rect 2584 407 2585 411
rect 2602 409 2621 413
rect 2679 411 2683 445
rect 2665 407 2673 411
rect 2678 409 2683 411
rect 2678 407 2905 409
rect 2485 388 2488 396
rect 2412 385 2423 387
rect 2485 385 2499 388
rect 2412 384 2417 385
rect 2193 381 2417 384
rect 2421 381 2423 385
rect 2193 380 2423 381
rect 2523 379 2526 406
rect 2585 397 2588 407
rect 2679 406 2905 407
rect 2692 405 2905 406
rect 2891 397 2895 398
rect 2585 393 2895 397
rect 2538 385 2597 388
rect 2428 376 2526 379
rect 2625 385 2887 388
rect 2611 381 2615 384
rect 2611 378 2678 381
rect 2179 373 2244 376
rect 2116 372 2169 373
rect 2034 369 2169 372
rect 2034 363 2037 369
rect 2241 366 2244 373
rect 2428 371 2432 376
rect 1983 360 2048 363
rect 1950 344 1991 348
rect 1987 337 1991 344
rect 1940 305 1941 309
rect 1948 335 1951 336
rect 1948 332 1955 335
rect 1948 267 1951 332
rect 1991 333 2024 336
rect 2044 336 2047 360
rect 2101 357 2109 360
rect 2126 360 2211 363
rect 2215 360 2236 363
rect 2312 362 2377 365
rect 2101 353 2103 357
rect 2107 355 2109 357
rect 2107 353 2176 355
rect 2101 352 2176 353
rect 2101 351 2109 352
rect 2095 332 2128 335
rect 2108 328 2111 332
rect 2220 328 2223 334
rect 2108 325 2223 328
rect 2184 316 2185 319
rect 2182 268 2185 316
rect 2233 310 2236 360
rect 2373 359 2377 362
rect 2428 359 2431 371
rect 2674 368 2678 378
rect 2435 365 2455 367
rect 2435 364 2451 365
rect 2435 360 2436 364
rect 2440 361 2451 364
rect 2455 362 2540 365
rect 2639 365 2704 368
rect 2440 360 2455 361
rect 2435 359 2443 360
rect 2373 356 2431 359
rect 2277 334 2284 337
rect 2227 306 2261 310
rect 2221 305 2261 306
rect 1948 264 2042 267
rect 2052 265 2195 268
rect 1912 248 1917 264
rect 2039 260 2042 264
rect 2006 250 2014 251
rect 2006 248 2007 250
rect 1912 244 2007 248
rect 2012 244 2014 250
rect 2006 242 2014 244
rect 2190 234 2221 238
rect 2171 233 2195 234
rect 2128 230 2195 233
rect 2128 229 2131 230
rect 2072 226 2131 229
rect 1897 220 1898 224
rect 2072 217 2076 226
rect 1982 214 2076 217
rect 1947 186 1954 189
rect 1947 121 1950 186
rect 1990 187 2023 190
rect 2043 190 2046 214
rect 2125 214 2210 217
rect 2178 204 2184 205
rect 2178 200 2179 204
rect 2183 200 2184 204
rect 2178 198 2184 200
rect 2004 152 2007 187
rect 2094 186 2127 189
rect 2107 182 2110 186
rect 2219 182 2222 188
rect 2107 179 2222 182
rect 2183 170 2184 173
rect 2104 154 2107 170
rect 2004 148 2097 152
rect 2103 151 2170 154
rect 2092 135 2097 148
rect 2092 131 2165 135
rect 2181 122 2184 170
rect 2234 166 2237 305
rect 2246 295 2259 299
rect 2245 282 2266 286
rect 2277 269 2280 334
rect 2320 335 2353 338
rect 2373 338 2376 356
rect 2512 354 2670 357
rect 2338 286 2342 335
rect 2424 334 2457 337
rect 2437 330 2440 334
rect 2549 330 2552 336
rect 2437 327 2552 330
rect 2604 337 2611 340
rect 2513 318 2514 321
rect 2511 270 2514 318
rect 2554 308 2588 312
rect 2548 307 2588 308
rect 2564 279 2592 282
rect 2604 272 2607 337
rect 2647 338 2680 341
rect 2700 341 2703 365
rect 2782 365 2867 368
rect 2759 357 2833 359
rect 2759 356 2837 357
rect 2663 283 2667 338
rect 2751 337 2784 340
rect 2764 333 2767 337
rect 2876 333 2879 339
rect 2764 330 2879 333
rect 2672 296 2675 321
rect 2840 321 2841 324
rect 2689 284 2748 287
rect 2756 283 2760 321
rect 2838 273 2841 321
rect 2277 266 2371 269
rect 2381 267 2524 270
rect 2604 269 2698 272
rect 2708 270 2851 273
rect 2256 258 2267 262
rect 2368 262 2371 266
rect 2695 265 2698 269
rect 2666 258 2686 261
rect 2256 253 2260 258
rect 2666 256 2669 258
rect 2426 253 2669 256
rect 2683 257 2686 258
rect 2746 258 2794 261
rect 2683 253 2685 257
rect 2689 253 2690 256
rect 2254 251 2264 253
rect 2254 245 2256 251
rect 2261 245 2264 251
rect 2254 243 2264 245
rect 2426 237 2429 253
rect 2746 249 2749 258
rect 2677 247 2749 249
rect 2673 246 2749 247
rect 2755 240 2760 243
rect 2246 234 2429 237
rect 2455 236 2760 240
rect 2455 235 2578 236
rect 2456 219 2461 235
rect 2788 222 2791 258
rect 2833 245 2866 248
rect 2835 230 2839 245
rect 2311 216 2376 219
rect 2343 200 2346 216
rect 2276 188 2283 191
rect 2229 165 2259 166
rect 2229 160 2258 165
rect 2199 131 2219 135
rect 1947 118 2041 121
rect 2051 119 2194 122
rect 2038 114 2041 118
rect 1939 79 1947 80
rect 1939 73 1941 79
rect 1945 75 1947 79
rect 1945 73 1966 75
rect 1939 72 1966 73
rect 1939 71 1969 72
rect 1864 19 1875 21
rect 1864 13 1866 19
rect 1873 13 1875 19
rect 1864 12 1875 13
rect 2230 17 2236 160
rect 2257 135 2261 136
rect 2245 131 2261 135
rect 2257 110 2261 131
rect 2276 123 2279 188
rect 2319 189 2352 192
rect 2372 192 2375 216
rect 2454 216 2539 219
rect 2638 219 2703 222
rect 2506 208 2513 209
rect 2506 203 2507 208
rect 2512 203 2513 208
rect 2506 201 2513 203
rect 2508 199 2512 201
rect 2334 142 2337 189
rect 2423 188 2456 191
rect 2436 184 2439 188
rect 2548 184 2551 190
rect 2436 181 2551 184
rect 2603 191 2610 194
rect 2343 176 2346 177
rect 2512 172 2513 175
rect 2343 150 2346 172
rect 2334 138 2433 142
rect 2510 124 2513 172
rect 2552 162 2588 165
rect 2526 138 2585 143
rect 2603 126 2606 191
rect 2646 192 2679 195
rect 2699 195 2702 219
rect 2781 219 2866 222
rect 2666 156 2670 192
rect 2750 191 2783 194
rect 2763 187 2766 191
rect 2875 187 2878 193
rect 2763 184 2878 187
rect 2839 175 2840 178
rect 2650 152 2670 156
rect 2666 151 2670 152
rect 2624 140 2751 143
rect 2757 140 2758 143
rect 2624 139 2758 140
rect 2837 127 2840 175
rect 2276 120 2370 123
rect 2380 121 2523 124
rect 2603 123 2697 126
rect 2707 124 2850 127
rect 2367 116 2370 120
rect 2694 119 2697 123
rect 2646 115 2650 116
rect 2257 106 2334 110
rect 2331 102 2334 106
rect 2414 105 2416 110
rect 2414 102 2419 105
rect 2315 73 2319 98
rect 2331 98 2419 102
rect 2331 97 2334 98
rect 2646 66 2650 111
rect 2884 105 2887 385
rect 2421 63 2650 66
rect 2421 62 2646 63
rect 2883 53 2887 105
rect 2388 49 2422 53
rect 2477 50 2887 53
rect 2883 49 2887 50
rect 2418 45 2422 49
rect 2418 42 2487 45
rect 2484 38 2487 42
rect 2891 38 2895 393
rect 2298 36 2301 38
rect 2292 32 2380 36
rect 2385 32 2465 35
rect 2484 34 2895 38
rect 2230 10 2231 17
rect 1496 4 1700 5
rect 1716 4 1832 5
rect 1496 3 1832 4
rect 1654 1 1832 3
rect 1580 -10 1582 -4
rect 1586 -8 1878 -4
rect 2298 -4 2301 32
rect 2902 24 2905 405
rect 2311 21 2905 24
rect 1586 -10 1881 -8
rect 2298 -9 2301 -8
<< metal3 >>
rect 1808 995 1906 997
rect 1808 994 1895 995
rect 1808 989 1812 994
rect 1817 991 1895 994
rect 1899 991 1906 995
rect 1817 989 1906 991
rect 1808 982 1819 989
rect 540 962 565 964
rect 540 958 541 962
rect 545 958 565 962
rect 540 957 546 958
rect 559 943 565 958
rect 1819 963 1829 965
rect 1819 961 1895 963
rect 1819 960 1886 961
rect 1819 953 1820 960
rect 1825 955 1886 960
rect 1894 955 1895 961
rect 1825 953 1895 955
rect 1819 950 1829 953
rect 559 941 566 943
rect 559 937 560 941
rect 564 937 566 941
rect 559 936 566 937
rect 1476 892 1534 893
rect 1476 887 1478 892
rect 1483 887 1534 892
rect 1476 886 1534 887
rect 1527 870 1534 886
rect 1527 869 1565 870
rect 1527 864 1558 869
rect 1563 864 1565 869
rect 1557 863 1565 864
rect 1841 869 1854 871
rect 1841 861 1844 869
rect 1850 861 1854 869
rect 1841 858 1854 861
rect 1843 823 1854 858
rect 1843 822 1945 823
rect 1843 813 1934 822
rect 1942 813 1945 822
rect 1843 812 1945 813
rect 1199 713 1214 714
rect 1199 709 1202 713
rect 1206 709 1214 713
rect 1199 706 1214 709
rect 1208 630 1214 706
rect 2019 644 2029 645
rect 2019 640 2023 644
rect 2027 640 2029 644
rect 2019 636 2029 640
rect 2261 643 2267 644
rect 2261 639 2262 643
rect 2266 639 2267 643
rect 1208 624 1274 630
rect 1056 617 1063 618
rect 1056 612 1057 617
rect 1062 612 1063 617
rect 321 597 336 598
rect 0 596 336 597
rect 0 591 326 596
rect 1 480 7 591
rect 321 589 326 591
rect 332 589 336 596
rect 321 586 336 589
rect 1056 587 1063 612
rect 1056 581 1231 587
rect 1223 570 1229 581
rect 1221 565 1229 570
rect 1221 558 1222 565
rect 1228 558 1229 565
rect 1221 557 1229 558
rect 1268 543 1274 624
rect 1342 627 1349 628
rect 1342 622 1343 627
rect 1348 622 1349 627
rect 1342 621 1349 622
rect 1343 571 1349 621
rect 2022 589 2028 636
rect 2022 585 2023 589
rect 2027 585 2028 589
rect 2022 584 2028 585
rect 2261 581 2267 639
rect 2261 577 2262 581
rect 2266 577 2267 581
rect 2261 576 2267 577
rect 1343 567 1344 571
rect 1348 567 1349 571
rect 1343 566 1349 567
rect 1224 536 1277 543
rect 2181 542 2189 543
rect 2181 538 2182 542
rect 2186 538 2189 542
rect 1224 492 1231 536
rect 1268 535 1274 536
rect 2102 521 2110 522
rect 2102 517 2104 521
rect 2108 517 2110 521
rect 1785 506 1796 507
rect 1899 506 1909 507
rect 1785 502 1909 506
rect 1785 495 1786 502
rect 1791 495 1909 502
rect 1785 494 1796 495
rect 1224 490 1234 492
rect 1224 486 1225 490
rect 1229 486 1234 490
rect 1224 484 1234 486
rect 28 480 37 482
rect 1 479 37 480
rect 1 474 31 479
rect 35 474 37 479
rect 28 471 37 474
rect 564 480 574 481
rect 564 476 568 480
rect 572 476 574 480
rect 564 475 574 476
rect 564 469 570 475
rect 564 463 704 469
rect 551 456 576 458
rect 551 452 552 456
rect 556 452 576 456
rect 551 451 557 452
rect 570 437 576 452
rect 570 435 577 437
rect 570 431 571 435
rect 575 431 577 435
rect 570 430 577 431
rect 698 400 704 463
rect 698 395 699 400
rect 703 395 704 400
rect 698 393 704 395
rect 1224 346 1231 484
rect 1899 466 1909 495
rect 2102 486 2110 517
rect 1900 443 1908 466
rect 1900 442 1912 443
rect 1900 435 1904 442
rect 1909 435 1912 442
rect 1900 432 1912 435
rect 1542 367 1551 369
rect 1542 361 1544 367
rect 1550 361 1551 367
rect 1542 360 1551 361
rect 2103 360 2109 486
rect 2181 476 2189 538
rect 2180 473 2189 476
rect 2180 408 2187 473
rect 2566 436 2611 437
rect 2566 432 2606 436
rect 2610 432 2611 436
rect 2566 431 2611 432
rect 2178 405 2188 408
rect 2178 400 2180 405
rect 2184 400 2188 405
rect 2178 398 2188 400
rect 2416 385 2441 387
rect 2416 381 2417 385
rect 2421 381 2441 385
rect 2416 380 2422 381
rect 1222 345 1231 346
rect 1222 341 1223 345
rect 1227 341 1231 345
rect 1222 337 1231 341
rect 729 322 735 323
rect 729 318 730 322
rect 734 318 735 322
rect 729 264 735 318
rect 454 217 465 219
rect 454 211 459 217
rect 464 211 465 217
rect 454 210 465 211
rect 458 159 465 210
rect 728 208 735 264
rect 1048 252 1090 253
rect 1048 248 1084 252
rect 1089 248 1090 252
rect 1048 247 1090 248
rect 1048 226 1054 247
rect 993 224 1054 226
rect 993 220 995 224
rect 1000 220 1054 224
rect 993 218 1054 220
rect 728 183 734 208
rect 1224 205 1231 337
rect 1543 307 1550 360
rect 2101 357 2109 360
rect 2435 366 2441 381
rect 2435 364 2442 366
rect 2435 360 2436 364
rect 2440 360 2442 364
rect 2435 359 2442 360
rect 2101 353 2103 357
rect 2107 353 2109 357
rect 2101 351 2109 353
rect 1543 301 1544 307
rect 1549 301 1550 307
rect 1543 299 1550 301
rect 1639 284 1649 286
rect 1639 278 1640 284
rect 1646 281 1649 284
rect 2566 282 2573 431
rect 1890 281 2574 282
rect 1646 278 2574 281
rect 1639 275 2574 278
rect 2254 251 2264 253
rect 2006 250 2014 251
rect 2006 244 2007 250
rect 2012 244 2014 250
rect 2006 242 2014 244
rect 2254 245 2256 251
rect 2261 250 2264 251
rect 2261 249 2320 250
rect 2261 248 2426 249
rect 2506 248 2513 252
rect 2261 245 2513 248
rect 2039 242 2184 243
rect 2006 236 2184 242
rect 2254 241 2513 245
rect 2254 240 2320 241
rect 2006 235 2151 236
rect 1651 226 1658 228
rect 1651 220 1652 226
rect 1657 225 1658 226
rect 1657 224 1903 225
rect 1657 220 1898 224
rect 1902 220 1903 224
rect 1651 219 1903 220
rect 1651 218 1658 219
rect 1222 204 1232 205
rect 1222 200 1223 204
rect 1227 200 1232 204
rect 1222 199 1232 200
rect 2178 204 2184 236
rect 2178 200 2179 204
rect 2183 200 2184 204
rect 2506 208 2513 241
rect 2506 203 2507 208
rect 2512 203 2513 208
rect 2506 201 2513 203
rect 2178 198 2184 200
rect 760 186 769 188
rect 728 180 740 183
rect 728 176 730 180
rect 734 176 740 180
rect 760 180 762 186
rect 767 184 769 186
rect 956 185 967 189
rect 906 184 967 185
rect 767 183 967 184
rect 767 181 965 183
rect 767 180 962 181
rect 760 177 962 180
rect 728 175 740 176
rect 950 176 961 177
rect 950 170 952 176
rect 958 170 961 176
rect 950 168 961 170
rect 458 158 676 159
rect 458 154 647 158
rect 652 154 676 158
rect 458 153 676 154
rect 668 87 676 153
rect 668 83 669 87
rect 673 83 676 87
rect 668 82 676 83
rect 951 52 961 168
rect 1940 79 1947 80
rect 1940 73 1941 79
rect 1945 73 1947 79
rect 1940 55 1947 73
rect 1786 53 1947 55
rect 951 46 954 52
rect 959 46 961 52
rect 951 44 961 46
rect 1578 51 1588 53
rect 1578 44 1581 51
rect 1586 44 1588 51
rect 1786 49 1787 53
rect 1791 49 1947 53
rect 1578 42 1588 44
rect 1579 -3 1588 42
rect 1625 45 1766 49
rect 1786 48 1795 49
rect 1625 39 1627 45
rect 1633 43 1766 45
rect 1633 39 1637 43
rect 1625 37 1637 39
rect 1760 31 1766 43
rect 1643 30 1650 31
rect 1643 26 1645 30
rect 1649 26 1650 30
rect 1643 17 1650 26
rect 1760 27 1761 31
rect 1765 27 1766 31
rect 1760 25 1766 27
rect 1864 19 1875 21
rect 1864 17 1866 19
rect 1643 13 1866 17
rect 1873 13 1875 19
rect 1643 11 1875 13
rect 1864 10 1875 11
rect 1579 -10 1582 -3
rect 1586 -10 1588 -3
rect 1579 -14 1588 -10
<< ntransistor >>
rect 1744 1048 1753 1050
rect 1744 1041 1753 1043
rect 164 1009 166 1020
rect 171 1009 173 1020
rect 184 1009 186 1018
rect 251 1009 253 1020
rect 258 1009 260 1020
rect 271 1009 273 1018
rect 344 1009 346 1020
rect 351 1009 353 1020
rect 364 1009 366 1018
rect 584 1011 586 1020
rect 597 1011 599 1022
rect 604 1011 606 1022
rect 677 1011 679 1020
rect 690 1011 692 1022
rect 697 1011 699 1022
rect 764 1011 766 1020
rect 777 1011 779 1022
rect 784 1011 786 1022
rect 1741 1029 1747 1031
rect 1625 1020 1631 1022
rect 1619 1008 1628 1010
rect 1619 1001 1628 1003
rect 1085 976 1087 979
rect 1741 1002 1753 1004
rect 1741 995 1753 997
rect 1741 985 1750 987
rect 1157 975 1159 978
rect 1196 975 1198 981
rect 1217 975 1219 981
rect 1250 975 1252 981
rect 1271 975 1273 981
rect 1306 975 1308 981
rect 1327 975 1329 981
rect 1360 975 1362 981
rect 1381 975 1383 981
rect 1741 975 1750 977
rect 1736 959 1745 961
rect 86 897 88 903
rect 98 891 100 900
rect 105 891 107 900
rect 164 899 166 908
rect 180 894 182 903
rect 190 894 192 903
rect 200 891 202 903
rect 207 891 209 903
rect 248 899 250 908
rect 264 894 266 903
rect 274 894 276 903
rect 284 891 286 903
rect 291 891 293 903
rect 318 897 320 903
rect 330 891 332 900
rect 337 891 339 900
rect 415 899 417 905
rect 427 893 429 902
rect 434 893 436 902
rect 493 901 495 910
rect 509 896 511 905
rect 519 896 521 905
rect 529 893 531 905
rect 536 893 538 905
rect 577 901 579 910
rect 593 896 595 905
rect 603 896 605 905
rect 613 893 615 905
rect 620 893 622 905
rect 647 899 649 905
rect 742 902 744 908
rect 1161 953 1163 956
rect 1200 950 1202 956
rect 1221 950 1223 956
rect 1254 950 1256 956
rect 1275 950 1277 956
rect 1310 950 1312 956
rect 1331 950 1333 956
rect 1364 950 1366 956
rect 1385 950 1387 956
rect 1627 942 1636 944
rect 659 893 661 902
rect 666 893 668 902
rect 754 896 756 905
rect 761 896 763 905
rect 820 904 822 913
rect 836 899 838 908
rect 846 899 848 908
rect 856 896 858 908
rect 863 896 865 908
rect 904 904 906 913
rect 920 899 922 908
rect 930 899 932 908
rect 940 896 942 908
rect 947 896 949 908
rect 974 902 976 908
rect 1591 927 1597 929
rect 1591 917 1597 919
rect 1591 907 1597 909
rect 986 896 988 905
rect 993 896 995 905
rect 1622 926 1631 928
rect 1622 916 1631 918
rect 1741 918 1753 920
rect 1741 911 1753 913
rect 1619 906 1631 908
rect 1619 899 1631 901
rect 1741 901 1750 903
rect 1741 891 1750 893
rect 179 863 181 869
rect 189 863 191 869
rect 199 863 201 869
rect 508 865 510 871
rect 518 865 520 871
rect 528 865 530 871
rect 835 868 837 874
rect 845 868 847 874
rect 855 868 857 874
rect 1775 910 1781 912
rect 1775 900 1781 902
rect 1775 890 1781 892
rect 2458 877 2460 883
rect 2468 877 2470 883
rect 2478 877 2480 883
rect 1736 875 1745 877
rect 2685 870 2687 883
rect 2695 873 2697 883
rect 2705 876 2707 890
rect 2715 876 2717 890
rect 2735 870 2737 890
rect 2742 870 2744 890
rect 2753 870 2755 884
rect 2818 879 2820 885
rect 2828 879 2830 885
rect 2838 879 2840 885
rect 1627 858 1636 860
rect 1085 831 1087 834
rect 1426 838 1428 848
rect 1157 830 1159 833
rect 1196 830 1198 836
rect 1217 830 1219 836
rect 1250 830 1252 836
rect 1271 830 1273 836
rect 1306 830 1308 836
rect 1327 830 1329 836
rect 1360 830 1362 836
rect 1381 830 1383 836
rect 1438 834 1440 848
rect 2320 846 2322 855
rect 2327 846 2329 855
rect 1622 842 1631 844
rect 1622 832 1631 834
rect 2339 843 2341 849
rect 2366 843 2368 855
rect 2373 843 2375 855
rect 2383 843 2385 852
rect 2393 843 2395 852
rect 2409 838 2411 847
rect 2450 843 2452 855
rect 2457 843 2459 855
rect 2467 843 2469 852
rect 2477 843 2479 852
rect 2493 838 2495 847
rect 2552 846 2554 855
rect 2559 846 2561 855
rect 1619 822 1631 824
rect 85 751 87 757
rect 97 745 99 754
rect 104 745 106 754
rect 163 753 165 762
rect 179 748 181 757
rect 189 748 191 757
rect 199 745 201 757
rect 206 745 208 757
rect 247 753 249 762
rect 263 748 265 757
rect 273 748 275 757
rect 283 745 285 757
rect 290 745 292 757
rect 317 751 319 757
rect 329 745 331 754
rect 336 745 338 754
rect 414 753 416 759
rect 426 747 428 756
rect 433 747 435 756
rect 492 755 494 764
rect 508 750 510 759
rect 518 750 520 759
rect 528 747 530 759
rect 535 747 537 759
rect 576 755 578 764
rect 592 750 594 759
rect 602 750 604 759
rect 612 747 614 759
rect 619 747 621 759
rect 646 753 648 759
rect 741 756 743 762
rect 1161 808 1163 811
rect 1200 805 1202 811
rect 1221 805 1223 811
rect 1254 805 1256 811
rect 1275 805 1277 811
rect 1310 805 1312 811
rect 1331 805 1333 811
rect 1364 805 1366 811
rect 1385 805 1387 811
rect 1619 815 1631 817
rect 1427 799 1429 809
rect 1439 799 1441 813
rect 1744 816 1753 818
rect 1744 809 1753 811
rect 1741 797 1747 799
rect 1625 788 1631 790
rect 658 747 660 756
rect 665 747 667 756
rect 753 750 755 759
rect 760 750 762 759
rect 819 758 821 767
rect 835 753 837 762
rect 845 753 847 762
rect 855 750 857 762
rect 862 750 864 762
rect 903 758 905 767
rect 919 753 921 762
rect 929 753 931 762
rect 939 750 941 762
rect 946 750 948 762
rect 973 756 975 762
rect 985 750 987 759
rect 992 750 994 759
rect 2571 843 2573 849
rect 2680 848 2682 857
rect 2687 848 2689 857
rect 2699 845 2701 851
rect 2726 845 2728 857
rect 2733 845 2735 857
rect 2743 845 2745 854
rect 2753 845 2755 854
rect 2769 840 2771 849
rect 2810 845 2812 857
rect 2817 845 2819 857
rect 2827 845 2829 854
rect 2837 845 2839 854
rect 2853 840 2855 849
rect 2912 848 2914 857
rect 2919 848 2921 857
rect 2931 845 2933 851
rect 1619 776 1628 778
rect 1619 769 1628 771
rect 178 717 180 723
rect 188 717 190 723
rect 198 717 200 723
rect 507 719 509 725
rect 517 719 519 725
rect 527 719 529 725
rect 834 722 836 728
rect 844 722 846 728
rect 854 722 856 728
rect 1992 735 1994 741
rect 2004 729 2006 738
rect 2011 729 2013 738
rect 2070 737 2072 746
rect 2086 732 2088 741
rect 2096 732 2098 741
rect 2106 729 2108 741
rect 2113 729 2115 741
rect 2154 737 2156 746
rect 2170 732 2172 741
rect 2180 732 2182 741
rect 2190 729 2192 741
rect 2197 729 2199 741
rect 2224 735 2226 741
rect 2236 729 2238 738
rect 2243 729 2245 738
rect 2348 727 2350 733
rect 2360 721 2362 730
rect 2367 721 2369 730
rect 2426 729 2428 738
rect 2442 724 2444 733
rect 2452 724 2454 733
rect 1084 689 1086 692
rect 1426 698 1428 708
rect 1156 688 1158 691
rect 1195 688 1197 694
rect 1216 688 1218 694
rect 1249 688 1251 694
rect 1270 688 1272 694
rect 1305 688 1307 694
rect 1326 688 1328 694
rect 1359 688 1361 694
rect 1380 688 1382 694
rect 1438 694 1440 708
rect 1989 703 1991 717
rect 2000 697 2002 717
rect 2007 697 2009 717
rect 2027 697 2029 711
rect 2037 697 2039 711
rect 2047 704 2049 714
rect 2057 704 2059 717
rect 2462 721 2464 733
rect 2469 721 2471 733
rect 2510 729 2512 738
rect 2526 724 2528 733
rect 2536 724 2538 733
rect 2546 721 2548 733
rect 2553 721 2555 733
rect 2580 727 2582 733
rect 2592 721 2594 730
rect 2599 721 2601 730
rect 2708 729 2710 735
rect 2720 723 2722 732
rect 2727 723 2729 732
rect 2786 731 2788 740
rect 2802 726 2804 735
rect 2812 726 2814 735
rect 2822 723 2824 735
rect 2829 723 2831 735
rect 2870 731 2872 740
rect 2886 726 2888 735
rect 2896 726 2898 735
rect 2906 723 2908 735
rect 2913 723 2915 735
rect 2940 729 2942 735
rect 2952 723 2954 732
rect 2959 723 2961 732
rect 1746 688 1755 690
rect 2085 701 2087 707
rect 2095 701 2097 707
rect 2105 701 2107 707
rect 1746 681 1755 683
rect 1160 666 1162 669
rect 1199 663 1201 669
rect 1220 663 1222 669
rect 1253 663 1255 669
rect 1274 663 1276 669
rect 1309 663 1311 669
rect 1330 663 1332 669
rect 1363 663 1365 669
rect 1384 663 1386 669
rect 1743 669 1749 671
rect 1627 660 1633 662
rect 2441 693 2443 699
rect 2451 693 2453 699
rect 2461 693 2463 699
rect 2801 695 2803 701
rect 2811 695 2813 701
rect 2821 695 2823 701
rect 1621 648 1630 650
rect 1621 641 1630 643
rect 1743 642 1755 644
rect 1743 635 1755 637
rect 1743 625 1752 627
rect 1743 615 1752 617
rect 379 603 381 612
rect 392 601 394 612
rect 399 601 401 612
rect 472 603 474 612
rect 485 601 487 612
rect 492 601 494 612
rect 559 603 561 612
rect 572 601 574 612
rect 579 601 581 612
rect 1738 599 1747 601
rect 1629 582 1638 584
rect 1593 567 1599 569
rect 1593 557 1599 559
rect 1593 547 1599 549
rect 1624 566 1633 568
rect 1624 556 1633 558
rect 1743 558 1755 560
rect 1743 551 1755 553
rect 1621 546 1633 548
rect 1621 539 1633 541
rect 1743 541 1752 543
rect 1743 531 1752 533
rect 175 503 177 514
rect 182 503 184 514
rect 195 503 197 512
rect 262 503 264 514
rect 269 503 271 514
rect 282 503 284 512
rect 355 503 357 514
rect 362 503 364 514
rect 375 503 377 512
rect 595 505 597 514
rect 608 505 610 516
rect 615 505 617 516
rect 688 505 690 514
rect 701 505 703 516
rect 708 505 710 516
rect 1777 550 1783 552
rect 1777 540 1783 542
rect 1777 530 1783 532
rect 775 505 777 514
rect 788 505 790 516
rect 795 505 797 516
rect 1738 515 1747 517
rect 1629 498 1638 500
rect 1106 465 1108 468
rect 1624 482 1633 484
rect 1624 472 1633 474
rect 1178 464 1180 467
rect 1217 464 1219 470
rect 1238 464 1240 470
rect 1271 464 1273 470
rect 1292 464 1294 470
rect 1327 464 1329 470
rect 1348 464 1350 470
rect 1381 464 1383 470
rect 1402 464 1404 470
rect 1621 462 1633 464
rect 1621 455 1633 457
rect 97 391 99 397
rect 109 385 111 394
rect 116 385 118 394
rect 175 393 177 402
rect 191 388 193 397
rect 201 388 203 397
rect 211 385 213 397
rect 218 385 220 397
rect 259 393 261 402
rect 275 388 277 397
rect 285 388 287 397
rect 295 385 297 397
rect 302 385 304 397
rect 329 391 331 397
rect 341 385 343 394
rect 348 385 350 394
rect 426 393 428 399
rect 438 387 440 396
rect 445 387 447 396
rect 504 395 506 404
rect 520 390 522 399
rect 530 390 532 399
rect 540 387 542 399
rect 547 387 549 399
rect 588 395 590 404
rect 604 390 606 399
rect 614 390 616 399
rect 624 387 626 399
rect 631 387 633 399
rect 658 393 660 399
rect 753 396 755 402
rect 1746 456 1755 458
rect 1746 449 1755 451
rect 1182 442 1184 445
rect 1221 439 1223 445
rect 1242 439 1244 445
rect 1275 439 1277 445
rect 1296 439 1298 445
rect 1331 439 1333 445
rect 1352 439 1354 445
rect 1385 439 1387 445
rect 1406 439 1408 445
rect 1743 437 1749 439
rect 1627 428 1633 430
rect 2040 432 2042 443
rect 2047 432 2049 443
rect 2060 432 2062 441
rect 2127 432 2129 443
rect 2134 432 2136 443
rect 2147 432 2149 441
rect 2220 432 2222 443
rect 2227 432 2229 443
rect 2240 432 2242 441
rect 2460 434 2462 443
rect 2473 434 2475 445
rect 2480 434 2482 445
rect 2553 434 2555 443
rect 2566 434 2568 445
rect 2573 434 2575 445
rect 2640 434 2642 443
rect 2653 434 2655 445
rect 2660 434 2662 445
rect 670 387 672 396
rect 677 387 679 396
rect 765 390 767 399
rect 772 390 774 399
rect 831 398 833 407
rect 847 393 849 402
rect 857 393 859 402
rect 867 390 869 402
rect 874 390 876 402
rect 915 398 917 407
rect 931 393 933 402
rect 941 393 943 402
rect 951 390 953 402
rect 958 390 960 402
rect 985 396 987 402
rect 1621 416 1630 418
rect 1621 409 1630 411
rect 997 390 999 399
rect 1004 390 1006 399
rect 190 357 192 363
rect 200 357 202 363
rect 210 357 212 363
rect 519 359 521 365
rect 529 359 531 365
rect 539 359 541 365
rect 846 362 848 368
rect 856 362 858 368
rect 866 362 868 368
rect 1104 320 1106 323
rect 1458 326 1460 336
rect 1470 326 1472 340
rect 1738 332 1747 334
rect 1176 319 1178 322
rect 1215 319 1217 325
rect 1236 319 1238 325
rect 1269 319 1271 325
rect 1290 319 1292 325
rect 1325 319 1327 325
rect 1346 319 1348 325
rect 1379 319 1381 325
rect 1400 319 1402 325
rect 1738 325 1747 327
rect 96 245 98 251
rect 108 239 110 248
rect 115 239 117 248
rect 174 247 176 256
rect 190 242 192 251
rect 200 242 202 251
rect 210 239 212 251
rect 217 239 219 251
rect 258 247 260 256
rect 274 242 276 251
rect 284 242 286 251
rect 294 239 296 251
rect 301 239 303 251
rect 328 245 330 251
rect 340 239 342 248
rect 347 239 349 248
rect 425 247 427 253
rect 437 241 439 250
rect 444 241 446 250
rect 503 249 505 258
rect 519 244 521 253
rect 529 244 531 253
rect 539 241 541 253
rect 546 241 548 253
rect 587 249 589 258
rect 603 244 605 253
rect 613 244 615 253
rect 623 241 625 253
rect 630 241 632 253
rect 657 247 659 253
rect 752 250 754 256
rect 1180 297 1182 300
rect 1219 294 1221 300
rect 1240 294 1242 300
rect 1273 294 1275 300
rect 1294 294 1296 300
rect 1329 294 1331 300
rect 1350 294 1352 300
rect 1383 294 1385 300
rect 1404 294 1406 300
rect 1962 320 1964 326
rect 1735 313 1741 315
rect 1974 314 1976 323
rect 1981 314 1983 323
rect 2040 322 2042 331
rect 2056 317 2058 326
rect 2066 317 2068 326
rect 2076 314 2078 326
rect 2083 314 2085 326
rect 2124 322 2126 331
rect 2140 317 2142 326
rect 2150 317 2152 326
rect 2160 314 2162 326
rect 2167 314 2169 326
rect 2194 320 2196 326
rect 2206 314 2208 323
rect 2213 314 2215 323
rect 2291 322 2293 328
rect 2303 316 2305 325
rect 2310 316 2312 325
rect 2369 324 2371 333
rect 2385 319 2387 328
rect 2395 319 2397 328
rect 2405 316 2407 328
rect 2412 316 2414 328
rect 2453 324 2455 333
rect 2469 319 2471 328
rect 2479 319 2481 328
rect 2489 316 2491 328
rect 2496 316 2498 328
rect 2523 322 2525 328
rect 2618 325 2620 331
rect 2535 316 2537 325
rect 2542 316 2544 325
rect 2630 319 2632 328
rect 2637 319 2639 328
rect 2696 327 2698 336
rect 2712 322 2714 331
rect 2722 322 2724 331
rect 2732 319 2734 331
rect 2739 319 2741 331
rect 2780 327 2782 336
rect 2796 322 2798 331
rect 2806 322 2808 331
rect 2816 319 2818 331
rect 2823 319 2825 331
rect 2850 325 2852 331
rect 2862 319 2864 328
rect 2869 319 2871 328
rect 1735 286 1747 288
rect 2055 286 2057 292
rect 2065 286 2067 292
rect 2075 286 2077 292
rect 2384 288 2386 294
rect 2394 288 2396 294
rect 2404 288 2406 294
rect 2711 291 2713 297
rect 2721 291 2723 297
rect 2731 291 2733 297
rect 1735 279 1747 281
rect 669 241 671 250
rect 676 241 678 250
rect 764 244 766 253
rect 771 244 773 253
rect 830 252 832 261
rect 846 247 848 256
rect 856 247 858 256
rect 866 244 868 256
rect 873 244 875 256
rect 914 252 916 261
rect 930 247 932 256
rect 940 247 942 256
rect 950 244 952 256
rect 957 244 959 256
rect 984 250 986 256
rect 1735 269 1744 271
rect 1735 259 1744 261
rect 996 244 998 253
rect 1003 244 1005 253
rect 189 211 191 217
rect 199 211 201 217
rect 209 211 211 217
rect 518 213 520 219
rect 528 213 530 219
rect 538 213 540 219
rect 845 216 847 222
rect 855 216 857 222
rect 865 216 867 222
rect 1730 243 1739 245
rect 1460 203 1462 213
rect 1472 199 1474 213
rect 1105 178 1107 181
rect 1735 202 1747 204
rect 1735 195 1747 197
rect 1735 185 1744 187
rect 1177 177 1179 180
rect 1216 177 1218 183
rect 1237 177 1239 183
rect 1270 177 1272 183
rect 1291 177 1293 183
rect 1326 177 1328 183
rect 1347 177 1349 183
rect 1380 177 1382 183
rect 1401 177 1403 183
rect 1735 175 1744 177
rect 1181 155 1183 158
rect 1220 152 1222 158
rect 1241 152 1243 158
rect 1274 152 1276 158
rect 1295 152 1297 158
rect 1330 152 1332 158
rect 1351 152 1353 158
rect 1384 152 1386 158
rect 1405 152 1407 158
rect 1462 147 1464 157
rect 1474 147 1476 161
rect 1769 194 1775 196
rect 1769 184 1775 186
rect 1769 174 1775 176
rect 1961 174 1963 180
rect 1973 168 1975 177
rect 1980 168 1982 177
rect 2039 176 2041 185
rect 2055 171 2057 180
rect 2065 171 2067 180
rect 2075 168 2077 180
rect 2082 168 2084 180
rect 2123 176 2125 185
rect 2139 171 2141 180
rect 2149 171 2151 180
rect 2159 168 2161 180
rect 2166 168 2168 180
rect 2193 174 2195 180
rect 2205 168 2207 177
rect 2212 168 2214 177
rect 2290 176 2292 182
rect 2302 170 2304 179
rect 2309 170 2311 179
rect 2368 178 2370 187
rect 2384 173 2386 182
rect 2394 173 2396 182
rect 2404 170 2406 182
rect 2411 170 2413 182
rect 2452 178 2454 187
rect 2468 173 2470 182
rect 2478 173 2480 182
rect 2488 170 2490 182
rect 2495 170 2497 182
rect 2522 176 2524 182
rect 2617 179 2619 185
rect 2534 170 2536 179
rect 2541 170 2543 179
rect 2629 173 2631 182
rect 2636 173 2638 182
rect 2695 181 2697 190
rect 2711 176 2713 185
rect 2721 176 2723 185
rect 2731 173 2733 185
rect 2738 173 2740 185
rect 2779 181 2781 190
rect 2795 176 2797 185
rect 2805 176 2807 185
rect 2815 173 2817 185
rect 2822 173 2824 185
rect 2849 179 2851 185
rect 2861 173 2863 182
rect 2868 173 2870 182
rect 1730 159 1739 161
rect 1759 146 1772 148
rect 1762 136 1772 138
rect 390 97 392 106
rect 403 95 405 106
rect 410 95 412 106
rect 483 97 485 106
rect 496 95 498 106
rect 503 95 505 106
rect 570 97 572 106
rect 583 95 585 106
rect 590 95 592 106
rect 2054 140 2056 146
rect 2064 140 2066 146
rect 2074 140 2076 146
rect 2383 142 2385 148
rect 2393 142 2395 148
rect 2403 142 2405 148
rect 2710 145 2712 151
rect 2720 145 2722 151
rect 2730 145 2732 151
rect 1765 126 1779 128
rect 1765 116 1779 118
rect 1738 100 1747 102
rect 1759 96 1779 98
rect 1738 93 1747 95
rect 1759 89 1779 91
rect 1735 81 1741 83
rect 1759 78 1773 80
rect 2255 26 2257 35
rect 2268 24 2270 35
rect 2275 24 2277 35
rect 2348 26 2350 35
rect 2361 24 2363 35
rect 2368 24 2370 35
rect 2435 26 2437 35
rect 2448 24 2450 35
rect 2455 24 2457 35
<< ptransistor >>
rect 1714 1049 1724 1051
rect 1714 1039 1724 1041
rect 1085 1012 1087 1018
rect 1712 1029 1724 1031
rect 1157 1012 1159 1018
rect 1196 1012 1198 1018
rect 1217 1012 1219 1018
rect 1250 1012 1252 1018
rect 1271 1012 1273 1018
rect 1306 1012 1308 1018
rect 1327 1012 1329 1018
rect 1360 1012 1362 1018
rect 1381 1012 1383 1018
rect 1648 1020 1660 1022
rect 164 974 166 987
rect 174 974 176 987
rect 184 976 186 994
rect 251 974 253 987
rect 261 974 263 987
rect 271 976 273 994
rect 344 974 346 987
rect 354 974 356 987
rect 364 976 366 994
rect 584 978 586 996
rect 594 976 596 989
rect 604 976 606 989
rect 677 978 679 996
rect 687 976 689 989
rect 697 976 699 989
rect 764 978 766 996
rect 1648 1010 1658 1012
rect 774 976 776 989
rect 784 976 786 989
rect 1648 1000 1658 1002
rect 1696 1003 1723 1005
rect 1705 993 1723 995
rect 1705 983 1723 985
rect 1696 967 1723 969
rect 86 920 88 932
rect 96 920 98 930
rect 106 920 108 930
rect 172 921 174 948
rect 188 921 190 939
rect 198 921 200 939
rect 208 921 210 948
rect 256 921 258 948
rect 272 921 274 939
rect 282 921 284 939
rect 292 921 294 948
rect 318 920 320 932
rect 328 920 330 930
rect 338 920 340 930
rect 415 922 417 934
rect 425 922 427 932
rect 435 922 437 932
rect 501 923 503 950
rect 517 923 519 941
rect 527 923 529 941
rect 537 923 539 950
rect 585 923 587 950
rect 601 923 603 941
rect 611 923 613 941
rect 621 923 623 950
rect 647 922 649 934
rect 657 922 659 932
rect 667 922 669 932
rect 742 925 744 937
rect 752 925 754 935
rect 762 925 764 935
rect 828 926 830 953
rect 844 926 846 944
rect 854 926 856 944
rect 864 926 866 953
rect 912 926 914 953
rect 928 926 930 944
rect 938 926 940 944
rect 948 926 950 953
rect 974 925 976 937
rect 984 925 986 935
rect 994 925 996 935
rect 1546 927 1564 929
rect 1546 920 1564 922
rect 1161 913 1163 919
rect 1200 913 1202 919
rect 1221 913 1223 919
rect 1254 913 1256 919
rect 1275 913 1277 919
rect 1310 913 1312 919
rect 1331 913 1333 919
rect 1364 913 1366 919
rect 1385 913 1387 919
rect 1555 907 1567 909
rect 1649 934 1676 936
rect 1649 918 1667 920
rect 1696 919 1723 921
rect 1649 908 1667 910
rect 1705 909 1723 911
rect 1649 898 1676 900
rect 1705 899 1723 901
rect 179 818 181 836
rect 186 818 188 836
rect 199 827 201 839
rect 1085 867 1087 873
rect 1157 867 1159 873
rect 1196 867 1198 873
rect 1217 867 1219 873
rect 1250 867 1252 873
rect 1271 867 1273 873
rect 1306 867 1308 873
rect 1327 867 1329 873
rect 1360 867 1362 873
rect 1381 867 1383 873
rect 1426 860 1428 877
rect 1438 860 1440 888
rect 1696 883 1723 885
rect 1805 910 1817 912
rect 2458 907 2460 919
rect 2471 910 2473 928
rect 2478 910 2480 928
rect 1808 897 1826 899
rect 2685 905 2687 930
rect 2698 905 2700 918
rect 1808 890 1826 892
rect 2708 902 2710 927
rect 2715 902 2717 927
rect 2733 902 2735 930
rect 2743 902 2745 930
rect 2753 902 2755 930
rect 2818 909 2820 921
rect 2831 912 2833 930
rect 2838 912 2840 930
rect 508 820 510 838
rect 515 820 517 838
rect 528 829 530 841
rect 835 823 837 841
rect 842 823 844 841
rect 855 832 857 844
rect 1649 850 1676 852
rect 1649 834 1667 836
rect 1649 824 1667 826
rect 85 774 87 786
rect 95 774 97 784
rect 105 774 107 784
rect 171 775 173 802
rect 187 775 189 793
rect 197 775 199 793
rect 207 775 209 802
rect 255 775 257 802
rect 271 775 273 793
rect 281 775 283 793
rect 291 775 293 802
rect 317 774 319 786
rect 327 774 329 784
rect 337 774 339 784
rect 414 776 416 788
rect 424 776 426 786
rect 434 776 436 786
rect 500 777 502 804
rect 516 777 518 795
rect 526 777 528 795
rect 536 777 538 804
rect 584 777 586 804
rect 600 777 602 795
rect 610 777 612 795
rect 620 777 622 804
rect 646 776 648 788
rect 656 776 658 786
rect 666 776 668 786
rect 741 779 743 791
rect 751 779 753 789
rect 761 779 763 789
rect 827 780 829 807
rect 843 780 845 798
rect 853 780 855 798
rect 863 780 865 807
rect 911 780 913 807
rect 927 780 929 798
rect 937 780 939 798
rect 947 780 949 807
rect 973 779 975 791
rect 1649 814 1676 816
rect 1714 817 1724 819
rect 2319 816 2321 826
rect 2329 816 2331 826
rect 2339 814 2341 826
rect 1714 807 1724 809
rect 1712 797 1724 799
rect 983 779 985 789
rect 993 779 995 789
rect 1161 768 1163 774
rect 1200 768 1202 774
rect 1221 768 1223 774
rect 1254 768 1256 774
rect 1275 768 1277 774
rect 1310 768 1312 774
rect 1331 768 1333 774
rect 1364 768 1366 774
rect 1385 768 1387 774
rect 1427 770 1429 787
rect 1439 759 1441 787
rect 1648 788 1660 790
rect 2365 798 2367 825
rect 2375 807 2377 825
rect 2385 807 2387 825
rect 2401 798 2403 825
rect 2449 798 2451 825
rect 2459 807 2461 825
rect 2469 807 2471 825
rect 2485 798 2487 825
rect 2551 816 2553 826
rect 2561 816 2563 826
rect 2571 814 2573 826
rect 2679 818 2681 828
rect 2689 818 2691 828
rect 2699 816 2701 828
rect 2725 800 2727 827
rect 2735 809 2737 827
rect 2745 809 2747 827
rect 2761 800 2763 827
rect 2809 800 2811 827
rect 2819 809 2821 827
rect 2829 809 2831 827
rect 2845 800 2847 827
rect 2911 818 2913 828
rect 2921 818 2923 828
rect 2931 816 2933 828
rect 1648 778 1658 780
rect 1648 768 1658 770
rect 1992 758 1994 770
rect 2002 758 2004 768
rect 2012 758 2014 768
rect 1084 725 1086 731
rect 1156 725 1158 731
rect 1195 725 1197 731
rect 1216 725 1218 731
rect 1249 725 1251 731
rect 1270 725 1272 731
rect 1305 725 1307 731
rect 1326 725 1328 731
rect 1359 725 1361 731
rect 1380 725 1382 731
rect 178 672 180 690
rect 185 672 187 690
rect 198 681 200 693
rect 1426 720 1428 737
rect 1438 720 1440 748
rect 2078 759 2080 786
rect 2094 759 2096 777
rect 2104 759 2106 777
rect 2114 759 2116 786
rect 2162 759 2164 786
rect 2178 759 2180 777
rect 2188 759 2190 777
rect 2198 759 2200 786
rect 2224 758 2226 770
rect 2234 758 2236 768
rect 2244 758 2246 768
rect 2348 750 2350 762
rect 2358 750 2360 760
rect 2368 750 2370 760
rect 2434 751 2436 778
rect 2450 751 2452 769
rect 2460 751 2462 769
rect 2470 751 2472 778
rect 2518 751 2520 778
rect 2534 751 2536 769
rect 2544 751 2546 769
rect 2554 751 2556 778
rect 2580 750 2582 762
rect 2590 750 2592 760
rect 2600 750 2602 760
rect 2708 752 2710 764
rect 2718 752 2720 762
rect 2728 752 2730 762
rect 507 674 509 692
rect 514 674 516 692
rect 527 683 529 695
rect 834 677 836 695
rect 841 677 843 695
rect 854 686 856 698
rect 1716 689 1726 691
rect 2794 753 2796 780
rect 2810 753 2812 771
rect 2820 753 2822 771
rect 2830 753 2832 780
rect 2878 753 2880 780
rect 2894 753 2896 771
rect 2904 753 2906 771
rect 2914 753 2916 780
rect 2940 752 2942 764
rect 2950 752 2952 762
rect 2960 752 2962 762
rect 1716 679 1726 681
rect 379 627 381 645
rect 389 634 391 647
rect 399 634 401 647
rect 472 627 474 645
rect 482 634 484 647
rect 492 634 494 647
rect 1714 669 1726 671
rect 1650 660 1662 662
rect 1989 657 1991 685
rect 1999 657 2001 685
rect 2009 657 2011 685
rect 2022 657 2024 685
rect 2027 657 2029 685
rect 2034 657 2036 685
rect 2044 669 2046 682
rect 2057 657 2059 682
rect 1650 650 1660 652
rect 559 627 561 645
rect 569 634 571 647
rect 579 634 581 647
rect 1650 640 1660 642
rect 1698 643 1725 645
rect 2085 656 2087 674
rect 2092 656 2094 674
rect 2105 665 2107 677
rect 2441 648 2443 666
rect 2448 648 2450 666
rect 2461 657 2463 669
rect 2801 650 2803 668
rect 2808 650 2810 668
rect 2821 659 2823 671
rect 1707 633 1725 635
rect 1160 626 1162 632
rect 1199 626 1201 632
rect 1220 626 1222 632
rect 1253 626 1255 632
rect 1274 626 1276 632
rect 1309 626 1311 632
rect 1330 626 1332 632
rect 1363 626 1365 632
rect 1384 626 1386 632
rect 1707 623 1725 625
rect 1698 607 1725 609
rect 1548 567 1566 569
rect 1548 560 1566 562
rect 1557 547 1569 549
rect 1651 574 1678 576
rect 1651 558 1669 560
rect 1698 559 1725 561
rect 1651 548 1669 550
rect 1707 549 1725 551
rect 1651 538 1678 540
rect 1707 539 1725 541
rect 1698 523 1725 525
rect 1807 550 1819 552
rect 1810 537 1828 539
rect 1810 530 1828 532
rect 175 468 177 481
rect 185 468 187 481
rect 195 470 197 488
rect 262 468 264 481
rect 272 468 274 481
rect 282 470 284 488
rect 355 468 357 481
rect 365 468 367 481
rect 375 470 377 488
rect 595 472 597 490
rect 605 470 607 483
rect 615 470 617 483
rect 688 472 690 490
rect 698 470 700 483
rect 708 470 710 483
rect 775 472 777 490
rect 1106 501 1108 507
rect 1178 501 1180 507
rect 1217 501 1219 507
rect 1238 501 1240 507
rect 1271 501 1273 507
rect 1292 501 1294 507
rect 1327 501 1329 507
rect 1348 501 1350 507
rect 1381 501 1383 507
rect 1402 501 1404 507
rect 785 470 787 483
rect 795 470 797 483
rect 1651 490 1678 492
rect 1651 474 1669 476
rect 1651 464 1669 466
rect 1651 454 1678 456
rect 97 414 99 426
rect 107 414 109 424
rect 117 414 119 424
rect 183 415 185 442
rect 199 415 201 433
rect 209 415 211 433
rect 219 415 221 442
rect 267 415 269 442
rect 283 415 285 433
rect 293 415 295 433
rect 303 415 305 442
rect 329 414 331 426
rect 339 414 341 424
rect 349 414 351 424
rect 426 416 428 428
rect 436 416 438 426
rect 446 416 448 426
rect 512 417 514 444
rect 528 417 530 435
rect 538 417 540 435
rect 548 417 550 444
rect 596 417 598 444
rect 612 417 614 435
rect 622 417 624 435
rect 632 417 634 444
rect 658 416 660 428
rect 668 416 670 426
rect 678 416 680 426
rect 753 419 755 431
rect 763 419 765 429
rect 773 419 775 429
rect 839 420 841 447
rect 855 420 857 438
rect 865 420 867 438
rect 875 420 877 447
rect 923 420 925 447
rect 939 420 941 438
rect 949 420 951 438
rect 959 420 961 447
rect 1716 457 1726 459
rect 1716 447 1726 449
rect 985 419 987 431
rect 995 419 997 429
rect 1005 419 1007 429
rect 1714 437 1726 439
rect 1650 428 1662 430
rect 1650 418 1660 420
rect 1182 402 1184 408
rect 1221 402 1223 408
rect 1242 402 1244 408
rect 1275 402 1277 408
rect 1296 402 1298 408
rect 1331 402 1333 408
rect 1352 402 1354 408
rect 1385 402 1387 408
rect 1406 402 1408 408
rect 1650 408 1660 410
rect 2040 397 2042 410
rect 2050 397 2052 410
rect 2060 399 2062 417
rect 2127 397 2129 410
rect 2137 397 2139 410
rect 2147 399 2149 417
rect 2220 397 2222 410
rect 2230 397 2232 410
rect 2240 399 2242 417
rect 2460 401 2462 419
rect 2470 399 2472 412
rect 2480 399 2482 412
rect 2553 401 2555 419
rect 2563 399 2565 412
rect 2573 399 2575 412
rect 2640 401 2642 419
rect 2650 399 2652 412
rect 2660 399 2662 412
rect 190 312 192 330
rect 197 312 199 330
rect 210 321 212 333
rect 1104 356 1106 362
rect 1176 356 1178 362
rect 1215 356 1217 362
rect 1236 356 1238 362
rect 1269 356 1271 362
rect 1290 356 1292 362
rect 1325 356 1327 362
rect 1346 356 1348 362
rect 1379 356 1381 362
rect 1400 356 1402 362
rect 519 314 521 332
rect 526 314 528 332
rect 539 323 541 335
rect 846 317 848 335
rect 853 317 855 335
rect 866 326 868 338
rect 1962 343 1964 355
rect 1972 343 1974 353
rect 1982 343 1984 353
rect 1708 333 1718 335
rect 1708 323 1718 325
rect 96 268 98 280
rect 106 268 108 278
rect 116 268 118 278
rect 182 269 184 296
rect 198 269 200 287
rect 208 269 210 287
rect 218 269 220 296
rect 266 269 268 296
rect 282 269 284 287
rect 292 269 294 287
rect 302 269 304 296
rect 328 268 330 280
rect 338 268 340 278
rect 348 268 350 278
rect 425 270 427 282
rect 435 270 437 280
rect 445 270 447 280
rect 511 271 513 298
rect 527 271 529 289
rect 537 271 539 289
rect 547 271 549 298
rect 595 271 597 298
rect 611 271 613 289
rect 621 271 623 289
rect 631 271 633 298
rect 657 270 659 282
rect 667 270 669 280
rect 677 270 679 280
rect 752 273 754 285
rect 762 273 764 283
rect 772 273 774 283
rect 838 274 840 301
rect 854 274 856 292
rect 864 274 866 292
rect 874 274 876 301
rect 922 274 924 301
rect 938 274 940 292
rect 948 274 950 292
rect 958 274 960 301
rect 984 273 986 285
rect 994 273 996 283
rect 1004 273 1006 283
rect 1458 297 1460 314
rect 1470 286 1472 314
rect 1706 313 1718 315
rect 2048 344 2050 371
rect 2064 344 2066 362
rect 2074 344 2076 362
rect 2084 344 2086 371
rect 2132 344 2134 371
rect 2148 344 2150 362
rect 2158 344 2160 362
rect 2168 344 2170 371
rect 2194 343 2196 355
rect 2204 343 2206 353
rect 2214 343 2216 353
rect 2291 345 2293 357
rect 2301 345 2303 355
rect 2311 345 2313 355
rect 2377 346 2379 373
rect 2393 346 2395 364
rect 2403 346 2405 364
rect 2413 346 2415 373
rect 2461 346 2463 373
rect 2477 346 2479 364
rect 2487 346 2489 364
rect 2497 346 2499 373
rect 2523 345 2525 357
rect 2533 345 2535 355
rect 2543 345 2545 355
rect 2618 348 2620 360
rect 2628 348 2630 358
rect 2638 348 2640 358
rect 2704 349 2706 376
rect 2720 349 2722 367
rect 2730 349 2732 367
rect 2740 349 2742 376
rect 2788 349 2790 376
rect 2804 349 2806 367
rect 2814 349 2816 367
rect 2824 349 2826 376
rect 2850 348 2852 360
rect 2860 348 2862 358
rect 2870 348 2872 358
rect 1690 287 1717 289
rect 1699 277 1717 279
rect 1699 267 1717 269
rect 1180 257 1182 263
rect 1219 257 1221 263
rect 1240 257 1242 263
rect 1273 257 1275 263
rect 1294 257 1296 263
rect 1329 257 1331 263
rect 1350 257 1352 263
rect 1383 257 1385 263
rect 1404 257 1406 263
rect 189 166 191 184
rect 196 166 198 184
rect 209 175 211 187
rect 1105 214 1107 220
rect 1460 225 1462 242
rect 1472 225 1474 253
rect 1690 251 1717 253
rect 2055 241 2057 259
rect 2062 241 2064 259
rect 2075 250 2077 262
rect 2384 243 2386 261
rect 2391 243 2393 261
rect 2404 252 2406 264
rect 2711 246 2713 264
rect 2718 246 2720 264
rect 2731 255 2733 267
rect 1177 214 1179 220
rect 1216 214 1218 220
rect 1237 214 1239 220
rect 1270 214 1272 220
rect 1291 214 1293 220
rect 1326 214 1328 220
rect 1347 214 1349 220
rect 1380 214 1382 220
rect 1401 214 1403 220
rect 518 168 520 186
rect 525 168 527 186
rect 538 177 540 189
rect 845 171 847 189
rect 852 171 854 189
rect 865 180 867 192
rect 1690 203 1717 205
rect 1699 193 1717 195
rect 1699 183 1717 185
rect 1690 167 1717 169
rect 390 121 392 139
rect 400 128 402 141
rect 410 128 412 141
rect 483 121 485 139
rect 493 128 495 141
rect 503 128 505 141
rect 570 121 572 139
rect 580 128 582 141
rect 590 128 592 141
rect 1961 197 1963 209
rect 1971 197 1973 207
rect 1981 197 1983 207
rect 1799 194 1811 196
rect 1802 181 1820 183
rect 1802 174 1820 176
rect 2047 198 2049 225
rect 2063 198 2065 216
rect 2073 198 2075 216
rect 2083 198 2085 225
rect 2131 198 2133 225
rect 2147 198 2149 216
rect 2157 198 2159 216
rect 2167 198 2169 225
rect 2193 197 2195 209
rect 2203 197 2205 207
rect 2213 197 2215 207
rect 2290 199 2292 211
rect 2300 199 2302 209
rect 2310 199 2312 209
rect 2376 200 2378 227
rect 2392 200 2394 218
rect 2402 200 2404 218
rect 2412 200 2414 227
rect 2460 200 2462 227
rect 2476 200 2478 218
rect 2486 200 2488 218
rect 2496 200 2498 227
rect 2522 199 2524 211
rect 2532 199 2534 209
rect 2542 199 2544 209
rect 2617 202 2619 214
rect 2627 202 2629 212
rect 2637 202 2639 212
rect 2703 203 2705 230
rect 2719 203 2721 221
rect 2729 203 2731 221
rect 2739 203 2741 230
rect 2787 203 2789 230
rect 2803 203 2805 221
rect 2813 203 2815 221
rect 2823 203 2825 230
rect 2849 202 2851 214
rect 2859 202 2861 212
rect 2869 202 2871 212
rect 1794 146 1819 148
rect 1181 115 1183 121
rect 1220 115 1222 121
rect 1241 115 1243 121
rect 1274 115 1276 121
rect 1295 115 1297 121
rect 1330 115 1332 121
rect 1351 115 1353 121
rect 1384 115 1386 121
rect 1405 115 1407 121
rect 1462 118 1464 135
rect 1474 107 1476 135
rect 1794 133 1807 135
rect 1791 123 1816 125
rect 1791 116 1816 118
rect 1708 101 1718 103
rect 1791 98 1819 100
rect 1708 91 1718 93
rect 2054 95 2056 113
rect 2061 95 2063 113
rect 2074 104 2076 116
rect 2383 97 2385 115
rect 2390 97 2392 115
rect 2403 106 2405 118
rect 2710 100 2712 118
rect 2717 100 2719 118
rect 2730 109 2732 121
rect 1706 81 1718 83
rect 1791 88 1819 90
rect 1791 78 1819 80
rect 2255 50 2257 68
rect 2265 57 2267 70
rect 2275 57 2277 70
rect 2348 50 2350 68
rect 2358 57 2360 70
rect 2368 57 2370 70
rect 2435 50 2437 68
rect 2445 57 2447 70
rect 2455 57 2457 70
<< polycontact >>
rect 1736 1049 1740 1053
rect 1704 1040 1708 1044
rect 1728 1030 1732 1034
rect 1640 1017 1644 1021
rect 171 999 175 1003
rect 181 999 185 1003
rect 161 991 165 995
rect 258 999 262 1003
rect 268 999 272 1003
rect 248 991 252 995
rect 351 999 355 1003
rect 361 999 365 1003
rect 341 991 345 995
rect 585 1001 589 1005
rect 595 1001 599 1005
rect 678 1001 682 1005
rect 688 1001 692 1005
rect 605 993 609 997
rect 765 1001 769 1005
rect 775 1001 779 1005
rect 698 993 702 997
rect 1083 997 1087 1001
rect 1664 1007 1668 1011
rect 785 993 789 997
rect 1155 996 1159 1000
rect 1193 996 1197 1000
rect 1214 996 1218 1000
rect 1247 996 1251 1000
rect 1268 996 1272 1000
rect 1303 996 1307 1000
rect 1324 996 1328 1000
rect 1357 996 1361 1000
rect 1378 996 1382 1000
rect 1632 998 1636 1002
rect 1727 1000 1731 1004
rect 1727 990 1731 994
rect 1733 969 1737 973
rect 97 936 101 940
rect 158 928 162 932
rect 87 912 91 916
rect 242 928 246 932
rect 195 913 199 917
rect 205 913 209 917
rect 329 936 333 940
rect 426 938 430 942
rect 487 930 491 934
rect 106 904 110 908
rect 174 907 178 911
rect 279 913 283 917
rect 289 913 293 917
rect 319 912 323 916
rect 258 907 262 911
rect 416 914 420 918
rect 338 904 342 908
rect 571 930 575 934
rect 524 915 528 919
rect 534 915 538 919
rect 658 938 662 942
rect 753 941 757 945
rect 814 933 818 937
rect 435 906 439 910
rect 503 909 507 913
rect 608 915 612 919
rect 618 915 622 919
rect 648 914 652 918
rect 587 909 591 913
rect 743 917 747 921
rect 667 906 671 910
rect 898 933 902 937
rect 851 918 855 922
rect 861 918 865 922
rect 985 941 989 945
rect 1712 953 1716 957
rect 1656 946 1660 950
rect 2708 947 2712 951
rect 1159 931 1163 935
rect 1197 931 1201 935
rect 1218 931 1222 935
rect 1251 931 1255 935
rect 1272 931 1276 935
rect 1307 931 1311 935
rect 1328 931 1332 935
rect 1361 931 1365 935
rect 1382 931 1386 935
rect 762 909 766 913
rect 830 912 834 916
rect 935 918 939 922
rect 945 918 949 922
rect 975 917 979 921
rect 914 912 918 916
rect 1578 928 1582 932
rect 1570 918 1574 922
rect 1578 916 1582 920
rect 994 909 998 913
rect 1577 908 1581 912
rect 1635 930 1639 934
rect 1641 909 1645 913
rect 1727 916 1731 920
rect 1641 899 1645 903
rect 1727 906 1731 910
rect 176 850 180 854
rect 188 850 192 854
rect 196 849 200 853
rect 505 852 509 856
rect 517 852 521 856
rect 186 842 190 846
rect 525 851 529 855
rect 832 855 836 859
rect 844 855 848 859
rect 515 844 519 848
rect 852 854 856 858
rect 842 847 846 851
rect 1083 852 1087 856
rect 1733 885 1737 889
rect 1791 907 1795 911
rect 1790 899 1794 903
rect 1798 897 1802 901
rect 2469 900 2473 904
rect 2459 893 2463 897
rect 2467 892 2471 896
rect 2479 892 2483 896
rect 1790 887 1794 891
rect 2692 897 2696 901
rect 2686 887 2690 891
rect 2706 894 2710 898
rect 2829 902 2833 906
rect 2725 894 2729 898
rect 2732 894 2736 898
rect 2742 894 2746 898
rect 2752 894 2756 898
rect 2819 895 2823 899
rect 2827 894 2831 898
rect 2839 894 2843 898
rect 1712 869 1716 873
rect 1656 862 1660 866
rect 1155 851 1159 855
rect 1193 851 1197 855
rect 1214 851 1218 855
rect 1247 851 1251 855
rect 1268 851 1272 855
rect 1303 851 1307 855
rect 1324 851 1328 855
rect 1357 851 1361 855
rect 1378 851 1382 855
rect 1423 852 1427 856
rect 1435 852 1439 856
rect 1635 846 1639 850
rect 2317 838 2321 842
rect 1641 825 1645 829
rect 2397 835 2401 839
rect 2336 830 2340 834
rect 2366 829 2370 833
rect 2376 829 2380 833
rect 2481 835 2485 839
rect 2549 838 2553 842
rect 96 790 100 794
rect 157 782 161 786
rect 86 766 90 770
rect 241 782 245 786
rect 194 767 198 771
rect 204 767 208 771
rect 328 790 332 794
rect 425 792 429 796
rect 486 784 490 788
rect 105 758 109 762
rect 173 761 177 765
rect 278 767 282 771
rect 288 767 292 771
rect 318 766 322 770
rect 257 761 261 765
rect 415 768 419 772
rect 337 758 341 762
rect 570 784 574 788
rect 523 769 527 773
rect 533 769 537 773
rect 657 792 661 796
rect 752 795 756 799
rect 813 787 817 791
rect 434 760 438 764
rect 502 763 506 767
rect 607 769 611 773
rect 617 769 621 773
rect 647 768 651 772
rect 586 763 590 767
rect 742 771 746 775
rect 666 760 670 764
rect 897 787 901 791
rect 850 772 854 776
rect 860 772 864 776
rect 984 795 988 799
rect 1641 815 1645 819
rect 1736 817 1740 821
rect 1704 808 1708 812
rect 1424 791 1428 795
rect 1436 791 1440 795
rect 1728 798 1732 802
rect 2326 806 2330 810
rect 1159 786 1163 790
rect 1197 786 1201 790
rect 1218 786 1222 790
rect 1251 786 1255 790
rect 1272 786 1276 790
rect 1307 786 1311 790
rect 1328 786 1332 790
rect 1361 786 1365 790
rect 1382 786 1386 790
rect 761 763 765 767
rect 829 766 833 770
rect 934 772 938 776
rect 944 772 948 776
rect 974 771 978 775
rect 913 766 917 770
rect 993 763 997 767
rect 1640 785 1644 789
rect 2450 829 2454 833
rect 2460 829 2464 833
rect 2413 814 2417 818
rect 2677 840 2681 844
rect 2568 830 2572 834
rect 2757 837 2761 841
rect 2696 832 2700 836
rect 2726 831 2730 835
rect 2736 831 2740 835
rect 2841 837 2845 841
rect 2909 840 2913 844
rect 2497 814 2501 818
rect 2558 806 2562 810
rect 2686 808 2690 812
rect 2810 831 2814 835
rect 2820 831 2824 835
rect 2773 816 2777 820
rect 2928 832 2932 836
rect 2857 816 2861 820
rect 2918 808 2922 812
rect 1664 775 1668 779
rect 1632 766 1636 770
rect 2003 774 2007 778
rect 2064 766 2068 770
rect 1993 750 1997 754
rect 175 704 179 708
rect 187 704 191 708
rect 195 703 199 707
rect 504 706 508 710
rect 516 706 520 710
rect 185 696 189 700
rect 524 705 528 709
rect 831 709 835 713
rect 843 709 847 713
rect 514 698 518 702
rect 851 708 855 712
rect 1082 710 1086 714
rect 2148 766 2152 770
rect 2101 751 2105 755
rect 2111 751 2115 755
rect 2235 774 2239 778
rect 2359 766 2363 770
rect 2012 742 2016 746
rect 2080 745 2084 749
rect 2185 751 2189 755
rect 2195 751 2199 755
rect 2225 750 2229 754
rect 2164 745 2168 749
rect 2420 758 2424 762
rect 2244 742 2248 746
rect 2349 742 2353 746
rect 2504 758 2508 762
rect 2457 743 2461 747
rect 2467 743 2471 747
rect 2591 766 2595 770
rect 2719 768 2723 772
rect 2780 760 2784 764
rect 2368 734 2372 738
rect 2436 737 2440 741
rect 2541 743 2545 747
rect 2551 743 2555 747
rect 2581 742 2585 746
rect 841 701 845 705
rect 1154 709 1158 713
rect 1192 709 1196 713
rect 1213 709 1217 713
rect 1246 709 1250 713
rect 1267 709 1271 713
rect 1302 709 1306 713
rect 1323 709 1327 713
rect 1356 709 1360 713
rect 1377 709 1381 713
rect 1423 712 1427 716
rect 1435 712 1439 716
rect 1738 689 1742 693
rect 2520 737 2524 741
rect 2709 744 2713 748
rect 2600 734 2604 738
rect 2864 760 2868 764
rect 2817 745 2821 749
rect 2827 745 2831 749
rect 2951 768 2955 772
rect 2728 736 2732 740
rect 2796 739 2800 743
rect 2901 745 2905 749
rect 2911 745 2915 749
rect 2941 744 2945 748
rect 2880 739 2884 743
rect 2960 736 2964 740
rect 1988 689 1992 693
rect 1998 689 2002 693
rect 2008 689 2012 693
rect 2015 689 2019 693
rect 2034 689 2038 693
rect 2054 696 2058 700
rect 1706 680 1710 684
rect 2048 686 2052 690
rect 400 626 404 630
rect 1730 670 1734 674
rect 1642 657 1646 661
rect 2082 688 2086 692
rect 2094 688 2098 692
rect 2102 687 2106 691
rect 2092 680 2096 684
rect 2438 680 2442 684
rect 2450 680 2454 684
rect 380 618 384 622
rect 390 618 394 622
rect 493 626 497 630
rect 1158 644 1162 648
rect 1196 644 1200 648
rect 1217 644 1221 648
rect 1250 644 1254 648
rect 1271 644 1275 648
rect 1306 644 1310 648
rect 1327 644 1331 648
rect 1360 644 1364 648
rect 1381 644 1385 648
rect 473 618 477 622
rect 483 618 487 622
rect 1666 647 1670 651
rect 1634 638 1638 642
rect 1729 640 1733 644
rect 2009 635 2013 639
rect 2458 679 2462 683
rect 2798 682 2802 686
rect 2810 682 2814 686
rect 2448 672 2452 676
rect 2818 681 2822 685
rect 2808 674 2812 678
rect 580 626 584 630
rect 1729 630 1733 634
rect 2033 633 2037 637
rect 560 618 564 622
rect 570 618 574 622
rect 1735 609 1739 613
rect 1714 593 1718 597
rect 1658 586 1662 590
rect 1580 568 1584 572
rect 1572 558 1576 562
rect 1580 556 1584 560
rect 1579 548 1583 552
rect 1637 570 1641 574
rect 1643 549 1647 553
rect 1729 556 1733 560
rect 1643 539 1647 543
rect 1729 546 1733 550
rect 1735 525 1739 529
rect 1793 547 1797 551
rect 1792 539 1796 543
rect 1800 537 1804 541
rect 1792 527 1796 531
rect 182 493 186 497
rect 192 493 196 497
rect 172 485 176 489
rect 269 493 273 497
rect 279 493 283 497
rect 259 485 263 489
rect 362 493 366 497
rect 372 493 376 497
rect 352 485 356 489
rect 596 495 600 499
rect 606 495 610 499
rect 689 495 693 499
rect 699 495 703 499
rect 616 487 620 491
rect 776 495 780 499
rect 786 495 790 499
rect 709 487 713 491
rect 1714 509 1718 513
rect 796 487 800 491
rect 1104 486 1108 490
rect 1658 502 1662 506
rect 1176 485 1180 489
rect 1214 485 1218 489
rect 1235 485 1239 489
rect 1268 485 1272 489
rect 1289 485 1293 489
rect 1324 485 1328 489
rect 1345 485 1349 489
rect 1378 485 1382 489
rect 1399 485 1403 489
rect 1637 486 1641 490
rect 1643 465 1647 469
rect 1643 455 1647 459
rect 108 430 112 434
rect 169 422 173 426
rect 98 406 102 410
rect 253 422 257 426
rect 206 407 210 411
rect 216 407 220 411
rect 340 430 344 434
rect 437 432 441 436
rect 498 424 502 428
rect 117 398 121 402
rect 185 401 189 405
rect 290 407 294 411
rect 300 407 304 411
rect 330 406 334 410
rect 269 401 273 405
rect 427 408 431 412
rect 349 398 353 402
rect 582 424 586 428
rect 535 409 539 413
rect 545 409 549 413
rect 669 432 673 436
rect 764 435 768 439
rect 825 427 829 431
rect 446 400 450 404
rect 514 403 518 407
rect 619 409 623 413
rect 629 409 633 413
rect 659 408 663 412
rect 598 403 602 407
rect 754 411 758 415
rect 678 400 682 404
rect 909 427 913 431
rect 862 412 866 416
rect 872 412 876 416
rect 1738 457 1742 461
rect 1706 448 1710 452
rect 996 435 1000 439
rect 1730 438 1734 442
rect 1180 420 1184 424
rect 1218 420 1222 424
rect 1239 420 1243 424
rect 1272 420 1276 424
rect 1293 420 1297 424
rect 1328 420 1332 424
rect 1349 420 1353 424
rect 1382 420 1386 424
rect 1403 420 1407 424
rect 1642 425 1646 429
rect 773 403 777 407
rect 841 406 845 410
rect 946 412 950 416
rect 956 412 960 416
rect 986 411 990 415
rect 925 406 929 410
rect 1666 415 1670 419
rect 2047 422 2051 426
rect 2057 422 2061 426
rect 1005 403 1009 407
rect 1634 406 1638 410
rect 2037 414 2041 418
rect 2134 422 2138 426
rect 2144 422 2148 426
rect 2124 414 2128 418
rect 2227 422 2231 426
rect 2237 422 2241 426
rect 2217 414 2221 418
rect 2461 424 2465 428
rect 2471 424 2475 428
rect 2554 424 2558 428
rect 2564 424 2568 428
rect 2481 416 2485 420
rect 2641 424 2645 428
rect 2651 424 2655 428
rect 2574 416 2578 420
rect 2661 416 2665 420
rect 187 344 191 348
rect 199 344 203 348
rect 207 343 211 347
rect 516 346 520 350
rect 528 346 532 350
rect 197 336 201 340
rect 536 345 540 349
rect 843 349 847 353
rect 855 349 859 353
rect 526 338 530 342
rect 863 348 867 352
rect 853 341 857 345
rect 1102 341 1106 345
rect 1973 359 1977 363
rect 1174 340 1178 344
rect 1212 340 1216 344
rect 1233 340 1237 344
rect 1266 340 1270 344
rect 1287 340 1291 344
rect 1322 340 1326 344
rect 1343 340 1347 344
rect 1376 340 1380 344
rect 1397 340 1401 344
rect 2034 351 2038 355
rect 1730 333 1734 337
rect 1963 335 1967 339
rect 1455 318 1459 322
rect 1467 318 1471 322
rect 1698 324 1702 328
rect 107 284 111 288
rect 168 276 172 280
rect 97 260 101 264
rect 252 276 256 280
rect 205 261 209 265
rect 215 261 219 265
rect 339 284 343 288
rect 436 286 440 290
rect 497 278 501 282
rect 116 252 120 256
rect 184 255 188 259
rect 289 261 293 265
rect 299 261 303 265
rect 329 260 333 264
rect 268 255 272 259
rect 426 262 430 266
rect 348 252 352 256
rect 581 278 585 282
rect 534 263 538 267
rect 544 263 548 267
rect 668 286 672 290
rect 763 289 767 293
rect 824 281 828 285
rect 445 254 449 258
rect 513 257 517 261
rect 618 263 622 267
rect 628 263 632 267
rect 658 262 662 266
rect 597 257 601 261
rect 753 265 757 269
rect 677 254 681 258
rect 908 281 912 285
rect 861 266 865 270
rect 871 266 875 270
rect 995 289 999 293
rect 1722 314 1726 318
rect 2118 351 2122 355
rect 2071 336 2075 340
rect 2081 336 2085 340
rect 2205 359 2209 363
rect 2302 361 2306 365
rect 2363 353 2367 357
rect 1982 327 1986 331
rect 2050 330 2054 334
rect 2155 336 2159 340
rect 2165 336 2169 340
rect 2195 335 2199 339
rect 2134 330 2138 334
rect 2292 337 2296 341
rect 2214 327 2218 331
rect 2447 353 2451 357
rect 2400 338 2404 342
rect 2410 338 2414 342
rect 2534 361 2538 365
rect 2629 364 2633 368
rect 2690 356 2694 360
rect 2311 329 2315 333
rect 2379 332 2383 336
rect 2484 338 2488 342
rect 2494 338 2498 342
rect 2524 337 2528 341
rect 2463 332 2467 336
rect 2619 340 2623 344
rect 2543 329 2547 333
rect 2774 356 2778 360
rect 2727 341 2731 345
rect 2737 341 2741 345
rect 2861 364 2865 368
rect 2638 332 2642 336
rect 2706 335 2710 339
rect 2811 341 2815 345
rect 2821 341 2825 345
rect 2851 340 2855 344
rect 2790 335 2794 339
rect 2870 332 2874 336
rect 1721 284 1725 288
rect 1178 275 1182 279
rect 1216 275 1220 279
rect 1237 275 1241 279
rect 1270 275 1274 279
rect 1291 275 1295 279
rect 1326 275 1330 279
rect 1347 275 1351 279
rect 1380 275 1384 279
rect 1401 275 1405 279
rect 772 257 776 261
rect 840 260 844 264
rect 945 266 949 270
rect 955 266 959 270
rect 985 265 989 269
rect 924 260 928 264
rect 1721 274 1725 278
rect 2052 273 2056 277
rect 2064 273 2068 277
rect 1004 257 1008 261
rect 1727 253 1731 257
rect 186 198 190 202
rect 198 198 202 202
rect 206 197 210 201
rect 515 200 519 204
rect 527 200 531 204
rect 196 190 200 194
rect 535 199 539 203
rect 2072 272 2076 276
rect 2381 275 2385 279
rect 2393 275 2397 279
rect 2062 265 2066 269
rect 1706 237 1710 241
rect 2401 274 2405 278
rect 2708 278 2712 282
rect 2720 278 2724 282
rect 2391 267 2395 271
rect 2728 277 2732 281
rect 2718 270 2722 274
rect 1457 217 1461 221
rect 1469 217 1473 221
rect 842 203 846 207
rect 854 203 858 207
rect 525 192 529 196
rect 862 202 866 206
rect 852 195 856 199
rect 1103 199 1107 203
rect 1175 198 1179 202
rect 1213 198 1217 202
rect 1234 198 1238 202
rect 1267 198 1271 202
rect 1288 198 1292 202
rect 1323 198 1327 202
rect 1344 198 1348 202
rect 1377 198 1381 202
rect 1398 198 1402 202
rect 1972 213 1976 217
rect 1721 200 1725 204
rect 1721 190 1725 194
rect 1727 169 1731 173
rect 411 120 415 124
rect 391 112 395 116
rect 401 112 405 116
rect 504 120 508 124
rect 2033 205 2037 209
rect 1785 191 1789 195
rect 1784 183 1788 187
rect 1792 181 1796 185
rect 1962 189 1966 193
rect 1784 171 1788 175
rect 2117 205 2121 209
rect 2070 190 2074 194
rect 2080 190 2084 194
rect 2204 213 2208 217
rect 2301 215 2305 219
rect 2362 207 2366 211
rect 1981 181 1985 185
rect 2049 184 2053 188
rect 2154 190 2158 194
rect 2164 190 2168 194
rect 2194 189 2198 193
rect 2133 184 2137 188
rect 2291 191 2295 195
rect 2213 181 2217 185
rect 2446 207 2450 211
rect 2399 192 2403 196
rect 2409 192 2413 196
rect 2533 215 2537 219
rect 2628 218 2632 222
rect 2689 210 2693 214
rect 2310 183 2314 187
rect 2378 186 2382 190
rect 2483 192 2487 196
rect 2493 192 2497 196
rect 2523 191 2527 195
rect 2462 186 2466 190
rect 2618 194 2622 198
rect 2542 183 2546 187
rect 2773 210 2777 214
rect 2726 195 2730 199
rect 2736 195 2740 199
rect 2860 218 2864 222
rect 2637 186 2641 190
rect 2705 189 2709 193
rect 2810 195 2814 199
rect 2820 195 2824 199
rect 2850 194 2854 198
rect 2789 189 2793 193
rect 2869 186 2873 190
rect 1706 153 1710 157
rect 1459 139 1463 143
rect 1471 139 1475 143
rect 1776 143 1780 147
rect 1179 133 1183 137
rect 1217 133 1221 137
rect 1238 133 1242 137
rect 1271 133 1275 137
rect 1292 133 1296 137
rect 1327 133 1331 137
rect 1348 133 1352 137
rect 1381 133 1385 137
rect 1402 133 1406 137
rect 1786 137 1790 141
rect 484 112 488 116
rect 494 112 498 116
rect 591 120 595 124
rect 571 112 575 116
rect 581 112 585 116
rect 1783 123 1787 127
rect 2051 127 2055 131
rect 2063 127 2067 131
rect 1730 101 1734 105
rect 1783 104 1787 108
rect 1698 92 1702 96
rect 1783 97 1787 101
rect 2071 126 2075 130
rect 2380 129 2384 133
rect 2392 129 2396 133
rect 2061 119 2065 123
rect 2400 128 2404 132
rect 2707 132 2711 136
rect 2719 132 2723 136
rect 2390 121 2394 125
rect 2727 131 2731 135
rect 2717 124 2721 128
rect 1722 82 1726 86
rect 1783 87 1787 91
rect 1783 77 1787 81
rect 2276 49 2280 53
rect 2256 41 2260 45
rect 2266 41 2270 45
rect 2369 49 2373 53
rect 2349 41 2353 45
rect 2359 41 2363 45
rect 2456 49 2460 53
rect 2436 41 2440 45
rect 2446 41 2450 45
rect 1812 12 1816 16
<< ndcontact >>
rect 1745 1052 1749 1056
rect 177 1025 181 1029
rect 264 1025 268 1029
rect 158 1015 162 1019
rect 357 1025 361 1029
rect 188 1013 192 1017
rect 245 1015 249 1019
rect 589 1027 593 1031
rect 275 1013 279 1017
rect 338 1015 342 1019
rect 682 1027 686 1031
rect 368 1013 372 1017
rect 578 1015 582 1019
rect 608 1017 612 1021
rect 769 1027 773 1031
rect 671 1015 675 1019
rect 701 1017 705 1021
rect 758 1015 762 1019
rect 788 1017 792 1021
rect 1626 1024 1630 1028
rect 1754 1034 1758 1038
rect 1614 1013 1618 1017
rect 1742 1023 1746 1027
rect 1070 976 1074 980
rect 1104 976 1108 980
rect 1142 975 1146 979
rect 1623 995 1627 999
rect 1754 1007 1758 1011
rect 1744 989 1748 993
rect 1176 975 1180 979
rect 1188 976 1192 980
rect 1222 976 1226 980
rect 1242 976 1246 980
rect 1276 976 1280 980
rect 1298 976 1302 980
rect 1332 976 1336 980
rect 1352 976 1356 980
rect 1386 976 1390 980
rect 1742 979 1746 983
rect 1745 967 1749 971
rect 80 898 84 902
rect 158 903 162 907
rect 242 903 246 907
rect 109 895 113 899
rect 172 895 176 899
rect 184 898 188 902
rect 194 896 198 900
rect 91 886 95 890
rect 256 895 260 899
rect 268 898 272 902
rect 278 896 282 900
rect 212 886 216 890
rect 312 898 316 902
rect 409 900 413 904
rect 487 905 491 909
rect 341 895 345 899
rect 571 905 575 909
rect 438 897 442 901
rect 501 897 505 901
rect 513 900 517 904
rect 523 898 527 902
rect 296 886 300 890
rect 323 886 327 890
rect 420 888 424 892
rect 585 897 589 901
rect 597 900 601 904
rect 607 898 611 902
rect 541 888 545 892
rect 641 900 645 904
rect 736 903 740 907
rect 1146 952 1150 956
rect 1180 952 1184 956
rect 1192 951 1196 955
rect 1226 951 1230 955
rect 1246 951 1250 955
rect 1280 951 1284 955
rect 1302 951 1306 955
rect 1336 951 1340 955
rect 1356 951 1360 955
rect 1390 951 1394 955
rect 1737 953 1741 957
rect 1631 946 1635 950
rect 814 908 818 912
rect 670 897 674 901
rect 898 908 902 912
rect 765 900 769 904
rect 828 900 832 904
rect 840 903 844 907
rect 850 901 854 905
rect 625 888 629 892
rect 652 888 656 892
rect 747 891 751 895
rect 912 900 916 904
rect 924 903 928 907
rect 934 901 938 905
rect 868 891 872 895
rect 968 903 972 907
rect 1592 931 1596 935
rect 1592 921 1596 925
rect 1592 911 1596 915
rect 997 900 1001 904
rect 1592 901 1596 905
rect 1623 932 1627 936
rect 1626 920 1630 924
rect 1754 923 1758 927
rect 1624 910 1628 914
rect 1744 905 1748 909
rect 952 891 956 895
rect 979 891 983 895
rect 1614 892 1618 896
rect 1742 895 1746 899
rect 173 864 177 868
rect 183 864 187 868
rect 193 864 197 868
rect 203 864 207 868
rect 502 866 506 870
rect 512 866 516 870
rect 522 866 526 870
rect 532 866 536 870
rect 829 869 833 873
rect 839 869 843 873
rect 849 869 853 873
rect 859 869 863 873
rect 1745 883 1749 887
rect 1776 914 1780 918
rect 1776 904 1780 908
rect 1776 894 1780 898
rect 1776 884 1780 888
rect 2452 878 2456 882
rect 2462 878 2466 882
rect 2472 878 2476 882
rect 2482 878 2486 882
rect 2679 878 2683 882
rect 1737 869 1741 873
rect 2689 874 2693 878
rect 2699 877 2703 881
rect 2709 885 2713 889
rect 2719 885 2723 889
rect 2719 878 2723 882
rect 2729 878 2733 882
rect 1631 862 1635 866
rect 2746 871 2750 875
rect 2757 878 2761 882
rect 2812 880 2816 884
rect 2822 880 2826 884
rect 2832 880 2836 884
rect 2842 880 2846 884
rect 1070 831 1074 835
rect 1104 831 1108 835
rect 1142 830 1146 834
rect 1420 843 1424 847
rect 1176 830 1180 834
rect 1188 831 1192 835
rect 1222 831 1226 835
rect 1242 831 1246 835
rect 1276 831 1280 835
rect 1298 831 1302 835
rect 1332 831 1336 835
rect 1352 831 1356 835
rect 1386 831 1390 835
rect 1431 835 1435 839
rect 1442 843 1446 847
rect 1442 836 1446 840
rect 1623 848 1627 852
rect 2332 856 2336 860
rect 2359 856 2363 860
rect 2314 847 2318 851
rect 1626 836 1630 840
rect 1624 826 1628 830
rect 2343 844 2347 848
rect 2443 856 2447 860
rect 2377 846 2381 850
rect 2387 844 2391 848
rect 2399 847 2403 851
rect 2564 856 2568 860
rect 2692 858 2696 862
rect 2719 858 2723 862
rect 2461 846 2465 850
rect 2471 844 2475 848
rect 2483 847 2487 851
rect 2546 847 2550 851
rect 2413 839 2417 843
rect 2674 849 2678 853
rect 2497 839 2501 843
rect 79 752 83 756
rect 157 757 161 761
rect 241 757 245 761
rect 108 749 112 753
rect 171 749 175 753
rect 183 752 187 756
rect 193 750 197 754
rect 90 740 94 744
rect 255 749 259 753
rect 267 752 271 756
rect 277 750 281 754
rect 211 740 215 744
rect 311 752 315 756
rect 408 754 412 758
rect 486 759 490 763
rect 340 749 344 753
rect 570 759 574 763
rect 437 751 441 755
rect 500 751 504 755
rect 512 754 516 758
rect 522 752 526 756
rect 295 740 299 744
rect 322 740 326 744
rect 419 742 423 746
rect 584 751 588 755
rect 596 754 600 758
rect 606 752 610 756
rect 540 742 544 746
rect 640 754 644 758
rect 735 757 739 761
rect 1146 807 1150 811
rect 1180 807 1184 811
rect 1192 806 1196 810
rect 1226 806 1230 810
rect 1246 806 1250 810
rect 1280 806 1284 810
rect 1302 806 1306 810
rect 1336 806 1340 810
rect 1356 806 1360 810
rect 1390 806 1394 810
rect 1421 800 1425 804
rect 1432 808 1436 812
rect 1443 807 1447 811
rect 1614 808 1618 812
rect 1745 820 1749 824
rect 1443 800 1447 804
rect 1626 792 1630 796
rect 1754 802 1758 806
rect 813 762 817 766
rect 669 751 673 755
rect 897 762 901 766
rect 764 754 768 758
rect 827 754 831 758
rect 839 757 843 761
rect 849 755 853 759
rect 624 742 628 746
rect 651 742 655 746
rect 746 745 750 749
rect 911 754 915 758
rect 923 757 927 761
rect 933 755 937 759
rect 867 745 871 749
rect 967 757 971 761
rect 996 754 1000 758
rect 1614 781 1618 785
rect 1742 791 1746 795
rect 2575 844 2579 848
rect 2703 846 2707 850
rect 2803 858 2807 862
rect 2737 848 2741 852
rect 2747 846 2751 850
rect 2759 849 2763 853
rect 2924 858 2928 862
rect 2821 848 2825 852
rect 2831 846 2835 850
rect 2843 849 2847 853
rect 2906 849 2910 853
rect 2773 841 2777 845
rect 2857 841 2861 845
rect 2935 846 2939 850
rect 1623 763 1627 767
rect 951 745 955 749
rect 978 745 982 749
rect 172 718 176 722
rect 182 718 186 722
rect 192 718 196 722
rect 202 718 206 722
rect 501 720 505 724
rect 511 720 515 724
rect 521 720 525 724
rect 531 720 535 724
rect 828 723 832 727
rect 838 723 842 727
rect 848 723 852 727
rect 858 723 862 727
rect 1986 736 1990 740
rect 2064 741 2068 745
rect 2148 741 2152 745
rect 2015 733 2019 737
rect 2078 733 2082 737
rect 2090 736 2094 740
rect 2100 734 2104 738
rect 1997 724 2001 728
rect 2162 733 2166 737
rect 2174 736 2178 740
rect 2184 734 2188 738
rect 2118 724 2122 728
rect 2218 736 2222 740
rect 2247 733 2251 737
rect 2202 724 2206 728
rect 2229 724 2233 728
rect 2342 728 2346 732
rect 2420 733 2424 737
rect 2504 733 2508 737
rect 2371 725 2375 729
rect 2434 725 2438 729
rect 2446 728 2450 732
rect 2456 726 2460 730
rect 1069 689 1073 693
rect 1103 689 1107 693
rect 1141 688 1145 692
rect 1420 703 1424 707
rect 1175 688 1179 692
rect 1187 689 1191 693
rect 1221 689 1225 693
rect 1241 689 1245 693
rect 1275 689 1279 693
rect 1297 689 1301 693
rect 1331 689 1335 693
rect 1351 689 1355 693
rect 1431 695 1435 699
rect 1442 703 1446 707
rect 1983 705 1987 709
rect 1994 712 1998 716
rect 1442 696 1446 700
rect 1385 689 1389 693
rect 1747 692 1751 696
rect 2011 705 2015 709
rect 2021 705 2025 709
rect 2021 698 2025 702
rect 2031 698 2035 702
rect 2041 706 2045 710
rect 2051 709 2055 713
rect 2353 716 2357 720
rect 2518 725 2522 729
rect 2530 728 2534 732
rect 2540 726 2544 730
rect 2474 716 2478 720
rect 2574 728 2578 732
rect 2702 730 2706 734
rect 2780 735 2784 739
rect 2603 725 2607 729
rect 2864 735 2868 739
rect 2731 727 2735 731
rect 2794 727 2798 731
rect 2806 730 2810 734
rect 2816 728 2820 732
rect 2558 716 2562 720
rect 2585 716 2589 720
rect 2713 718 2717 722
rect 2878 727 2882 731
rect 2890 730 2894 734
rect 2900 728 2904 732
rect 2834 718 2838 722
rect 2934 730 2938 734
rect 2963 727 2967 731
rect 2918 718 2922 722
rect 2945 718 2949 722
rect 2061 705 2065 709
rect 2079 702 2083 706
rect 2089 702 2093 706
rect 2099 702 2103 706
rect 2109 702 2113 706
rect 1145 665 1149 669
rect 1179 665 1183 669
rect 1191 664 1195 668
rect 1225 664 1229 668
rect 1245 664 1249 668
rect 1279 664 1283 668
rect 1301 664 1305 668
rect 1335 664 1339 668
rect 1355 664 1359 668
rect 1389 664 1393 668
rect 1628 664 1632 668
rect 1756 674 1760 678
rect 1616 653 1620 657
rect 1744 663 1748 667
rect 2435 694 2439 698
rect 2445 694 2449 698
rect 2455 694 2459 698
rect 2465 694 2469 698
rect 2795 696 2799 700
rect 2805 696 2809 700
rect 2815 696 2819 700
rect 2825 696 2829 700
rect 1625 635 1629 639
rect 1756 647 1760 651
rect 1746 629 1750 633
rect 1744 619 1748 623
rect 373 604 377 608
rect 403 602 407 606
rect 466 604 470 608
rect 496 602 500 606
rect 553 604 557 608
rect 384 592 388 596
rect 583 602 587 606
rect 477 592 481 596
rect 1747 607 1751 611
rect 564 592 568 596
rect 1739 593 1743 597
rect 1633 586 1637 590
rect 1594 571 1598 575
rect 1594 561 1598 565
rect 1594 551 1598 555
rect 1594 541 1598 545
rect 1625 572 1629 576
rect 1628 560 1632 564
rect 1756 563 1760 567
rect 1626 550 1630 554
rect 1746 545 1750 549
rect 1616 532 1620 536
rect 1744 535 1748 539
rect 188 519 192 523
rect 275 519 279 523
rect 169 509 173 513
rect 368 519 372 523
rect 199 507 203 511
rect 256 509 260 513
rect 600 521 604 525
rect 286 507 290 511
rect 349 509 353 513
rect 693 521 697 525
rect 379 507 383 511
rect 589 509 593 513
rect 619 511 623 515
rect 780 521 784 525
rect 682 509 686 513
rect 712 511 716 515
rect 1747 523 1751 527
rect 1778 554 1782 558
rect 1778 544 1782 548
rect 1778 534 1782 538
rect 1778 524 1782 528
rect 769 509 773 513
rect 799 511 803 515
rect 1739 509 1743 513
rect 1633 502 1637 506
rect 1091 465 1095 469
rect 1125 465 1129 469
rect 1163 464 1167 468
rect 1625 488 1629 492
rect 1628 476 1632 480
rect 1197 464 1201 468
rect 1209 465 1213 469
rect 1243 465 1247 469
rect 1263 465 1267 469
rect 1297 465 1301 469
rect 1319 465 1323 469
rect 1353 465 1357 469
rect 1373 465 1377 469
rect 1407 465 1411 469
rect 1626 466 1630 470
rect 91 392 95 396
rect 169 397 173 401
rect 253 397 257 401
rect 120 389 124 393
rect 183 389 187 393
rect 195 392 199 396
rect 205 390 209 394
rect 102 380 106 384
rect 267 389 271 393
rect 279 392 283 396
rect 289 390 293 394
rect 223 380 227 384
rect 323 392 327 396
rect 420 394 424 398
rect 498 399 502 403
rect 352 389 356 393
rect 582 399 586 403
rect 449 391 453 395
rect 512 391 516 395
rect 524 394 528 398
rect 534 392 538 396
rect 307 380 311 384
rect 334 380 338 384
rect 431 382 435 386
rect 596 391 600 395
rect 608 394 612 398
rect 618 392 622 396
rect 552 382 556 386
rect 652 394 656 398
rect 747 397 751 401
rect 1616 448 1620 452
rect 1747 460 1751 464
rect 2053 448 2057 452
rect 1167 441 1171 445
rect 1201 441 1205 445
rect 1213 440 1217 444
rect 1247 440 1251 444
rect 1267 440 1271 444
rect 1301 440 1305 444
rect 1323 440 1327 444
rect 1357 440 1361 444
rect 1377 440 1381 444
rect 1411 440 1415 444
rect 1628 432 1632 436
rect 1756 442 1760 446
rect 2140 448 2144 452
rect 2034 438 2038 442
rect 1616 421 1620 425
rect 1744 431 1748 435
rect 2233 448 2237 452
rect 2064 436 2068 440
rect 2121 438 2125 442
rect 2465 450 2469 454
rect 2151 436 2155 440
rect 2214 438 2218 442
rect 2558 450 2562 454
rect 2244 436 2248 440
rect 2454 438 2458 442
rect 2484 440 2488 444
rect 2645 450 2649 454
rect 2547 438 2551 442
rect 2577 440 2581 444
rect 2634 438 2638 442
rect 2664 440 2668 444
rect 825 402 829 406
rect 681 391 685 395
rect 909 402 913 406
rect 776 394 780 398
rect 839 394 843 398
rect 851 397 855 401
rect 861 395 865 399
rect 636 382 640 386
rect 663 382 667 386
rect 758 385 762 389
rect 923 394 927 398
rect 935 397 939 401
rect 945 395 949 399
rect 879 385 883 389
rect 979 397 983 401
rect 1625 403 1629 407
rect 1008 394 1012 398
rect 963 385 967 389
rect 990 385 994 389
rect 184 358 188 362
rect 194 358 198 362
rect 204 358 208 362
rect 214 358 218 362
rect 513 360 517 364
rect 523 360 527 364
rect 533 360 537 364
rect 543 360 547 364
rect 840 363 844 367
rect 850 363 854 367
rect 860 363 864 367
rect 870 363 874 367
rect 1089 320 1093 324
rect 1123 320 1127 324
rect 1161 319 1165 323
rect 1452 327 1456 331
rect 1463 335 1467 339
rect 1474 334 1478 338
rect 1474 327 1478 331
rect 1739 336 1743 340
rect 1195 319 1199 323
rect 1207 320 1211 324
rect 1241 320 1245 324
rect 1261 320 1265 324
rect 1295 320 1299 324
rect 1317 320 1321 324
rect 1351 320 1355 324
rect 1371 320 1375 324
rect 1405 320 1409 324
rect 90 246 94 250
rect 168 251 172 255
rect 252 251 256 255
rect 119 243 123 247
rect 182 243 186 247
rect 194 246 198 250
rect 204 244 208 248
rect 101 234 105 238
rect 266 243 270 247
rect 278 246 282 250
rect 288 244 292 248
rect 222 234 226 238
rect 322 246 326 250
rect 419 248 423 252
rect 497 253 501 257
rect 351 243 355 247
rect 581 253 585 257
rect 448 245 452 249
rect 511 245 515 249
rect 523 248 527 252
rect 533 246 537 250
rect 306 234 310 238
rect 333 234 337 238
rect 430 236 434 240
rect 595 245 599 249
rect 607 248 611 252
rect 617 246 621 250
rect 551 236 555 240
rect 651 248 655 252
rect 746 251 750 255
rect 1165 296 1169 300
rect 1199 296 1203 300
rect 1211 295 1215 299
rect 1245 295 1249 299
rect 1265 295 1269 299
rect 1299 295 1303 299
rect 1321 295 1325 299
rect 1355 295 1359 299
rect 1375 295 1379 299
rect 1409 295 1413 299
rect 1748 318 1752 322
rect 1956 321 1960 325
rect 2034 326 2038 330
rect 2118 326 2122 330
rect 1985 318 1989 322
rect 2048 318 2052 322
rect 2060 321 2064 325
rect 2070 319 2074 323
rect 1736 307 1740 311
rect 1967 309 1971 313
rect 2132 318 2136 322
rect 2144 321 2148 325
rect 2154 319 2158 323
rect 2088 309 2092 313
rect 2188 321 2192 325
rect 2285 323 2289 327
rect 2363 328 2367 332
rect 2217 318 2221 322
rect 2447 328 2451 332
rect 2314 320 2318 324
rect 2377 320 2381 324
rect 2389 323 2393 327
rect 2399 321 2403 325
rect 2172 309 2176 313
rect 2199 309 2203 313
rect 2296 311 2300 315
rect 2461 320 2465 324
rect 2473 323 2477 327
rect 2483 321 2487 325
rect 2417 311 2421 315
rect 2517 323 2521 327
rect 2612 326 2616 330
rect 2690 331 2694 335
rect 2546 320 2550 324
rect 2774 331 2778 335
rect 2641 323 2645 327
rect 2704 323 2708 327
rect 2716 326 2720 330
rect 2726 324 2730 328
rect 2501 311 2505 315
rect 2528 311 2532 315
rect 2623 314 2627 318
rect 2788 323 2792 327
rect 2800 326 2804 330
rect 2810 324 2814 328
rect 2744 314 2748 318
rect 2844 326 2848 330
rect 2873 323 2877 327
rect 2828 314 2832 318
rect 2855 314 2859 318
rect 1748 291 1752 295
rect 2049 287 2053 291
rect 2059 287 2063 291
rect 2069 287 2073 291
rect 2079 287 2083 291
rect 2378 289 2382 293
rect 2388 289 2392 293
rect 2398 289 2402 293
rect 2408 289 2412 293
rect 2705 292 2709 296
rect 2715 292 2719 296
rect 2725 292 2729 296
rect 2735 292 2739 296
rect 824 256 828 260
rect 680 245 684 249
rect 908 256 912 260
rect 775 248 779 252
rect 838 248 842 252
rect 850 251 854 255
rect 860 249 864 253
rect 635 236 639 240
rect 662 236 666 240
rect 757 239 761 243
rect 922 248 926 252
rect 934 251 938 255
rect 944 249 948 253
rect 878 239 882 243
rect 978 251 982 255
rect 1738 273 1742 277
rect 1736 263 1740 267
rect 1007 248 1011 252
rect 962 239 966 243
rect 989 239 993 243
rect 183 212 187 216
rect 193 212 197 216
rect 203 212 207 216
rect 213 212 217 216
rect 512 214 516 218
rect 522 214 526 218
rect 532 214 536 218
rect 542 214 546 218
rect 839 217 843 221
rect 849 217 853 221
rect 859 217 863 221
rect 869 217 873 221
rect 1739 251 1743 255
rect 1731 237 1735 241
rect 1454 208 1458 212
rect 1090 178 1094 182
rect 1465 200 1469 204
rect 1476 208 1480 212
rect 1748 207 1752 211
rect 1476 201 1480 205
rect 1124 178 1128 182
rect 1162 177 1166 181
rect 1738 189 1742 193
rect 1196 177 1200 181
rect 1208 178 1212 182
rect 1242 178 1246 182
rect 1262 178 1266 182
rect 1296 178 1300 182
rect 1318 178 1322 182
rect 1352 178 1356 182
rect 1372 178 1376 182
rect 1406 178 1410 182
rect 1736 179 1740 183
rect 1166 154 1170 158
rect 1200 154 1204 158
rect 1212 153 1216 157
rect 1246 153 1250 157
rect 1266 153 1270 157
rect 1300 153 1304 157
rect 1322 153 1326 157
rect 1356 153 1360 157
rect 1376 153 1380 157
rect 1410 153 1414 157
rect 1456 148 1460 152
rect 1467 156 1471 160
rect 1739 167 1743 171
rect 1770 198 1774 202
rect 1770 188 1774 192
rect 1770 178 1774 182
rect 1770 168 1774 172
rect 1955 175 1959 179
rect 2033 180 2037 184
rect 2117 180 2121 184
rect 1984 172 1988 176
rect 2047 172 2051 176
rect 2059 175 2063 179
rect 2069 173 2073 177
rect 1966 163 1970 167
rect 2131 172 2135 176
rect 2143 175 2147 179
rect 2153 173 2157 177
rect 2087 163 2091 167
rect 2187 175 2191 179
rect 2284 177 2288 181
rect 2362 182 2366 186
rect 2216 172 2220 176
rect 2446 182 2450 186
rect 2313 174 2317 178
rect 2376 174 2380 178
rect 2388 177 2392 181
rect 2398 175 2402 179
rect 2171 163 2175 167
rect 2198 163 2202 167
rect 2295 165 2299 169
rect 2460 174 2464 178
rect 2472 177 2476 181
rect 2482 175 2486 179
rect 2416 165 2420 169
rect 2516 177 2520 181
rect 2611 180 2615 184
rect 2689 185 2693 189
rect 2545 174 2549 178
rect 2773 185 2777 189
rect 2640 177 2644 181
rect 2703 177 2707 181
rect 2715 180 2719 184
rect 2725 178 2729 182
rect 2500 165 2504 169
rect 2527 165 2531 169
rect 2622 168 2626 172
rect 2787 177 2791 181
rect 2799 180 2803 184
rect 2809 178 2813 182
rect 2743 168 2747 172
rect 2843 180 2847 184
rect 2872 177 2876 181
rect 2827 168 2831 172
rect 2854 168 2858 172
rect 1478 155 1482 159
rect 1731 153 1735 157
rect 1478 148 1482 152
rect 1767 150 1771 154
rect 1763 140 1767 144
rect 384 98 388 102
rect 414 96 418 100
rect 477 98 481 102
rect 507 96 511 100
rect 564 98 568 102
rect 395 86 399 90
rect 1766 130 1770 134
rect 2048 141 2052 145
rect 2058 141 2062 145
rect 2068 141 2072 145
rect 2078 141 2082 145
rect 2377 143 2381 147
rect 2387 143 2391 147
rect 2397 143 2401 147
rect 2407 143 2411 147
rect 2704 146 2708 150
rect 2714 146 2718 150
rect 2724 146 2728 150
rect 2734 146 2738 150
rect 1774 120 1778 124
rect 1767 110 1771 114
rect 1774 110 1778 114
rect 594 96 598 100
rect 488 86 492 90
rect 1739 104 1743 108
rect 1767 100 1771 104
rect 575 86 579 90
rect 1748 86 1752 90
rect 1760 83 1764 87
rect 1736 75 1740 79
rect 1767 72 1771 76
rect 2249 27 2253 31
rect 2279 25 2283 29
rect 2342 27 2346 31
rect 2372 25 2376 29
rect 2429 27 2433 31
rect 2260 15 2264 19
rect 2459 25 2463 29
rect 2353 15 2357 19
rect 2440 15 2444 19
<< pdcontact >>
rect 1715 1053 1719 1057
rect 1719 1043 1723 1047
rect 1059 1013 1063 1017
rect 1103 1013 1109 1019
rect 1719 1033 1723 1037
rect 1649 1024 1653 1028
rect 1719 1023 1723 1027
rect 1142 1013 1146 1017
rect 1175 1013 1179 1017
rect 1188 1013 1192 1017
rect 1205 1013 1209 1017
rect 1222 1013 1226 1017
rect 1242 1013 1246 1017
rect 1259 1013 1263 1017
rect 1276 1013 1280 1017
rect 1298 1013 1302 1017
rect 1315 1013 1319 1017
rect 1332 1013 1336 1017
rect 1352 1013 1356 1017
rect 1369 1013 1373 1017
rect 1386 1013 1390 1017
rect 1649 1014 1653 1018
rect 158 975 162 979
rect 168 982 172 986
rect 168 975 172 979
rect 178 977 182 981
rect 188 989 192 993
rect 188 982 192 986
rect 245 975 249 979
rect 255 982 259 986
rect 255 975 259 979
rect 265 977 269 981
rect 275 989 279 993
rect 275 982 279 986
rect 338 975 342 979
rect 348 982 352 986
rect 348 975 352 979
rect 358 977 362 981
rect 368 989 372 993
rect 368 982 372 986
rect 578 991 582 995
rect 578 984 582 988
rect 671 991 675 995
rect 588 979 592 983
rect 598 984 602 988
rect 598 977 602 981
rect 671 984 675 988
rect 608 977 612 981
rect 758 991 762 995
rect 681 979 685 983
rect 691 984 695 988
rect 691 977 695 981
rect 758 984 762 988
rect 701 977 705 981
rect 1649 1004 1653 1008
rect 768 979 772 983
rect 778 984 782 988
rect 778 977 782 981
rect 788 977 792 981
rect 1653 994 1657 998
rect 1703 1007 1707 1011
rect 1711 997 1715 1001
rect 1718 987 1722 991
rect 1697 971 1701 975
rect 1704 971 1708 975
rect 1718 961 1722 965
rect 80 921 84 925
rect 90 921 94 925
rect 100 921 104 925
rect 110 925 114 929
rect 166 922 170 926
rect 176 943 180 947
rect 176 936 180 940
rect 192 922 196 926
rect 202 929 206 933
rect 212 937 216 941
rect 250 922 254 926
rect 260 943 264 947
rect 260 936 264 940
rect 276 922 280 926
rect 286 929 290 933
rect 296 937 300 941
rect 312 921 316 925
rect 322 921 326 925
rect 332 921 336 925
rect 342 925 346 929
rect 409 923 413 927
rect 419 923 423 927
rect 429 923 433 927
rect 439 927 443 931
rect 495 924 499 928
rect 505 945 509 949
rect 505 938 509 942
rect 521 924 525 928
rect 531 931 535 935
rect 541 939 545 943
rect 579 924 583 928
rect 589 945 593 949
rect 589 938 593 942
rect 605 924 609 928
rect 615 931 619 935
rect 625 939 629 943
rect 641 923 645 927
rect 651 923 655 927
rect 661 923 665 927
rect 671 927 675 931
rect 736 926 740 930
rect 746 926 750 930
rect 756 926 760 930
rect 766 930 770 934
rect 822 927 826 931
rect 832 948 836 952
rect 832 941 836 945
rect 848 927 852 931
rect 858 934 862 938
rect 868 942 872 946
rect 906 927 910 931
rect 916 948 920 952
rect 916 941 920 945
rect 932 927 936 931
rect 942 934 946 938
rect 952 942 956 946
rect 968 926 972 930
rect 978 926 982 930
rect 988 926 992 930
rect 998 930 1002 934
rect 1554 931 1558 935
rect 1146 914 1150 918
rect 1179 914 1183 918
rect 1192 914 1196 918
rect 1209 914 1213 918
rect 1226 914 1230 918
rect 1246 914 1250 918
rect 1263 914 1267 918
rect 1280 914 1284 918
rect 1302 914 1306 918
rect 1319 914 1323 918
rect 1336 914 1340 918
rect 1356 914 1360 918
rect 1373 914 1377 918
rect 1390 914 1394 918
rect 1547 913 1551 917
rect 1556 901 1560 905
rect 1650 938 1654 942
rect 1664 928 1668 932
rect 1671 928 1675 932
rect 1703 923 1707 927
rect 2464 923 2468 927
rect 1650 912 1654 916
rect 1711 913 1715 917
rect 1657 902 1661 906
rect 1718 903 1722 907
rect 1431 886 1435 890
rect 1665 892 1669 896
rect 1059 868 1063 872
rect 173 826 177 830
rect 1103 868 1109 874
rect 1142 868 1146 872
rect 1175 868 1179 872
rect 1188 868 1192 872
rect 1205 868 1209 872
rect 1222 868 1226 872
rect 1242 868 1246 872
rect 1259 868 1263 872
rect 1276 868 1280 872
rect 1298 868 1302 872
rect 1315 868 1319 872
rect 1332 868 1336 872
rect 1352 868 1356 872
rect 1369 868 1373 872
rect 1386 868 1390 872
rect 1420 868 1424 872
rect 1697 887 1701 891
rect 1704 887 1708 891
rect 1442 876 1446 880
rect 1718 877 1722 881
rect 1812 914 1816 918
rect 2452 914 2456 918
rect 2482 916 2486 920
rect 2679 913 2683 917
rect 1821 902 1825 906
rect 2679 906 2683 910
rect 2690 925 2694 929
rect 2702 906 2706 910
rect 1814 884 1818 888
rect 2725 925 2729 929
rect 2725 918 2729 922
rect 2737 917 2741 921
rect 2737 910 2741 914
rect 2747 925 2751 929
rect 2747 918 2751 922
rect 2824 925 2828 929
rect 2812 916 2816 920
rect 2757 910 2761 914
rect 2842 918 2846 922
rect 2757 903 2761 907
rect 1442 869 1446 873
rect 203 828 207 832
rect 502 828 506 832
rect 191 819 195 823
rect 532 830 536 834
rect 829 831 833 835
rect 520 821 524 825
rect 859 833 863 837
rect 1650 854 1654 858
rect 1664 844 1668 848
rect 1671 844 1675 848
rect 847 824 851 828
rect 1650 828 1654 832
rect 79 775 83 779
rect 89 775 93 779
rect 99 775 103 779
rect 109 779 113 783
rect 165 776 169 780
rect 175 797 179 801
rect 175 790 179 794
rect 191 776 195 780
rect 201 783 205 787
rect 211 791 215 795
rect 249 776 253 780
rect 259 797 263 801
rect 259 790 263 794
rect 275 776 279 780
rect 285 783 289 787
rect 295 791 299 795
rect 311 775 315 779
rect 321 775 325 779
rect 331 775 335 779
rect 341 779 345 783
rect 408 777 412 781
rect 418 777 422 781
rect 428 777 432 781
rect 438 781 442 785
rect 494 778 498 782
rect 504 799 508 803
rect 504 792 508 796
rect 520 778 524 782
rect 530 785 534 789
rect 540 793 544 797
rect 578 778 582 782
rect 588 799 592 803
rect 588 792 592 796
rect 604 778 608 782
rect 614 785 618 789
rect 624 793 628 797
rect 640 777 644 781
rect 650 777 654 781
rect 660 777 664 781
rect 670 781 674 785
rect 735 780 739 784
rect 745 780 749 784
rect 755 780 759 784
rect 765 784 769 788
rect 821 781 825 785
rect 831 802 835 806
rect 831 795 835 799
rect 847 781 851 785
rect 857 788 861 792
rect 867 796 871 800
rect 905 781 909 785
rect 915 802 919 806
rect 915 795 919 799
rect 931 781 935 785
rect 941 788 945 792
rect 951 796 955 800
rect 967 780 971 784
rect 1657 818 1661 822
rect 1665 808 1669 812
rect 1715 821 1719 825
rect 2313 817 2317 821
rect 2323 821 2327 825
rect 2333 821 2337 825
rect 1719 811 1723 815
rect 2343 821 2347 825
rect 1719 801 1723 805
rect 2359 805 2363 809
rect 1649 792 1653 796
rect 1719 791 1723 795
rect 977 780 981 784
rect 987 780 991 784
rect 997 784 1001 788
rect 1421 775 1425 779
rect 1146 769 1150 773
rect 1179 769 1183 773
rect 1192 769 1196 773
rect 1209 769 1213 773
rect 1226 769 1230 773
rect 1246 769 1250 773
rect 1263 769 1267 773
rect 1280 769 1284 773
rect 1302 769 1306 773
rect 1319 769 1323 773
rect 1336 769 1340 773
rect 1356 769 1360 773
rect 1373 769 1377 773
rect 1390 769 1394 773
rect 1432 757 1436 761
rect 1649 782 1653 786
rect 2369 813 2373 817
rect 2379 820 2383 824
rect 2395 806 2399 810
rect 2395 799 2399 803
rect 2405 820 2409 824
rect 2443 805 2447 809
rect 2453 813 2457 817
rect 2463 820 2467 824
rect 2479 806 2483 810
rect 2479 799 2483 803
rect 2489 820 2493 824
rect 2545 817 2549 821
rect 2555 821 2559 825
rect 2565 821 2569 825
rect 2575 821 2579 825
rect 2673 819 2677 823
rect 2683 823 2687 827
rect 2693 823 2697 827
rect 2703 823 2707 827
rect 2719 807 2723 811
rect 2729 815 2733 819
rect 2739 822 2743 826
rect 2755 808 2759 812
rect 2755 801 2759 805
rect 2765 822 2769 826
rect 2803 807 2807 811
rect 2813 815 2817 819
rect 2823 822 2827 826
rect 2839 808 2843 812
rect 2839 801 2843 805
rect 2849 822 2853 826
rect 2905 819 2909 823
rect 2915 823 2919 827
rect 2925 823 2929 827
rect 2935 823 2939 827
rect 1443 774 1447 778
rect 1649 772 1653 776
rect 1443 767 1447 771
rect 1653 762 1657 766
rect 1986 759 1990 763
rect 1996 759 2000 763
rect 2006 759 2010 763
rect 2016 763 2020 767
rect 1431 746 1435 750
rect 1058 726 1062 730
rect 1102 726 1108 732
rect 1141 726 1145 730
rect 1174 726 1178 730
rect 1187 726 1191 730
rect 1204 726 1208 730
rect 1221 726 1225 730
rect 1241 726 1245 730
rect 1258 726 1262 730
rect 1275 726 1279 730
rect 1297 726 1301 730
rect 1314 726 1318 730
rect 1331 726 1335 730
rect 1351 726 1355 730
rect 1368 726 1372 730
rect 1385 726 1389 730
rect 1420 728 1424 732
rect 172 680 176 684
rect 1442 736 1446 740
rect 2072 760 2076 764
rect 2082 781 2086 785
rect 2082 774 2086 778
rect 2098 760 2102 764
rect 2108 767 2112 771
rect 2118 775 2122 779
rect 2156 760 2160 764
rect 2166 781 2170 785
rect 2166 774 2170 778
rect 2182 760 2186 764
rect 2192 767 2196 771
rect 2202 775 2206 779
rect 2218 759 2222 763
rect 2228 759 2232 763
rect 2238 759 2242 763
rect 2248 763 2252 767
rect 1442 729 1446 733
rect 2342 751 2346 755
rect 2352 751 2356 755
rect 2362 751 2366 755
rect 2372 755 2376 759
rect 2428 752 2432 756
rect 2438 773 2442 777
rect 2438 766 2442 770
rect 2454 752 2458 756
rect 2464 759 2468 763
rect 2474 767 2478 771
rect 2512 752 2516 756
rect 2522 773 2526 777
rect 2522 766 2526 770
rect 2538 752 2542 756
rect 2548 759 2552 763
rect 2558 767 2562 771
rect 2574 751 2578 755
rect 2584 751 2588 755
rect 2594 751 2598 755
rect 2604 755 2608 759
rect 2702 753 2706 757
rect 2712 753 2716 757
rect 2722 753 2726 757
rect 2732 757 2736 761
rect 202 682 206 686
rect 501 682 505 686
rect 190 673 194 677
rect 531 684 535 688
rect 828 685 832 689
rect 519 675 523 679
rect 858 687 862 691
rect 1717 693 1721 697
rect 2788 754 2792 758
rect 2798 775 2802 779
rect 2798 768 2802 772
rect 2814 754 2818 758
rect 2824 761 2828 765
rect 2834 769 2838 773
rect 2872 754 2876 758
rect 2882 775 2886 779
rect 2882 768 2886 772
rect 2898 754 2902 758
rect 2908 761 2912 765
rect 2918 769 2922 773
rect 2934 753 2938 757
rect 2944 753 2948 757
rect 2954 753 2958 757
rect 2964 757 2968 761
rect 846 678 850 682
rect 1721 683 1725 687
rect 1983 680 1987 684
rect 373 635 377 639
rect 373 628 377 632
rect 383 640 387 644
rect 393 642 397 646
rect 393 635 397 639
rect 403 642 407 646
rect 466 635 470 639
rect 466 628 470 632
rect 476 640 480 644
rect 486 642 490 646
rect 486 635 490 639
rect 496 642 500 646
rect 1721 673 1725 677
rect 1983 673 1987 677
rect 1651 664 1655 668
rect 1721 663 1725 667
rect 1651 654 1655 658
rect 1993 665 1997 669
rect 1993 658 1997 662
rect 2003 673 2007 677
rect 2003 666 2007 670
rect 2015 665 2019 669
rect 2015 658 2019 662
rect 2038 677 2042 681
rect 2050 658 2054 662
rect 2061 677 2065 681
rect 2061 670 2065 674
rect 2079 664 2083 668
rect 553 635 557 639
rect 553 628 557 632
rect 563 640 567 644
rect 573 642 577 646
rect 573 635 577 639
rect 583 642 587 646
rect 1651 644 1655 648
rect 1655 634 1659 638
rect 1705 647 1709 651
rect 1713 637 1717 641
rect 2109 666 2113 670
rect 2097 657 2101 661
rect 2435 656 2439 660
rect 2465 658 2469 662
rect 2795 658 2799 662
rect 2453 649 2457 653
rect 2825 660 2829 664
rect 2813 651 2817 655
rect 1145 627 1149 631
rect 1178 627 1182 631
rect 1191 627 1195 631
rect 1208 627 1212 631
rect 1225 627 1229 631
rect 1245 627 1249 631
rect 1262 627 1266 631
rect 1279 627 1283 631
rect 1301 627 1305 631
rect 1318 627 1322 631
rect 1335 627 1339 631
rect 1355 627 1359 631
rect 1372 627 1376 631
rect 1389 627 1393 631
rect 1720 627 1724 631
rect 1699 611 1703 615
rect 1706 611 1710 615
rect 1720 601 1724 605
rect 1556 571 1560 575
rect 1549 553 1553 557
rect 1558 541 1562 545
rect 1652 578 1656 582
rect 1666 568 1670 572
rect 1673 568 1677 572
rect 1705 563 1709 567
rect 1652 552 1656 556
rect 1713 553 1717 557
rect 1659 542 1663 546
rect 1720 543 1724 547
rect 1667 532 1671 536
rect 1699 527 1703 531
rect 1706 527 1710 531
rect 1720 517 1724 521
rect 1814 554 1818 558
rect 1823 542 1827 546
rect 1816 524 1820 528
rect 169 469 173 473
rect 179 476 183 480
rect 179 469 183 473
rect 189 471 193 475
rect 199 483 203 487
rect 199 476 203 480
rect 256 469 260 473
rect 266 476 270 480
rect 266 469 270 473
rect 276 471 280 475
rect 286 483 290 487
rect 286 476 290 480
rect 349 469 353 473
rect 359 476 363 480
rect 359 469 363 473
rect 369 471 373 475
rect 379 483 383 487
rect 379 476 383 480
rect 589 485 593 489
rect 589 478 593 482
rect 682 485 686 489
rect 599 473 603 477
rect 609 478 613 482
rect 609 471 613 475
rect 682 478 686 482
rect 619 471 623 475
rect 769 485 773 489
rect 692 473 696 477
rect 702 478 706 482
rect 702 471 706 475
rect 769 478 773 482
rect 712 471 716 475
rect 1080 502 1084 506
rect 1124 502 1130 508
rect 1163 502 1167 506
rect 1196 502 1200 506
rect 1209 502 1213 506
rect 1226 502 1230 506
rect 1243 502 1247 506
rect 1263 502 1267 506
rect 1280 502 1284 506
rect 1297 502 1301 506
rect 1319 502 1323 506
rect 1336 502 1340 506
rect 1353 502 1357 506
rect 1373 502 1377 506
rect 1390 502 1394 506
rect 1407 502 1411 506
rect 779 473 783 477
rect 789 478 793 482
rect 789 471 793 475
rect 799 471 803 475
rect 1652 494 1656 498
rect 1666 484 1670 488
rect 1673 484 1677 488
rect 1652 468 1656 472
rect 1659 458 1663 462
rect 91 415 95 419
rect 101 415 105 419
rect 111 415 115 419
rect 121 419 125 423
rect 177 416 181 420
rect 187 437 191 441
rect 187 430 191 434
rect 203 416 207 420
rect 213 423 217 427
rect 223 431 227 435
rect 261 416 265 420
rect 271 437 275 441
rect 271 430 275 434
rect 287 416 291 420
rect 297 423 301 427
rect 307 431 311 435
rect 323 415 327 419
rect 333 415 337 419
rect 343 415 347 419
rect 353 419 357 423
rect 420 417 424 421
rect 430 417 434 421
rect 440 417 444 421
rect 450 421 454 425
rect 506 418 510 422
rect 516 439 520 443
rect 516 432 520 436
rect 532 418 536 422
rect 542 425 546 429
rect 552 433 556 437
rect 590 418 594 422
rect 600 439 604 443
rect 600 432 604 436
rect 616 418 620 422
rect 626 425 630 429
rect 636 433 640 437
rect 652 417 656 421
rect 662 417 666 421
rect 672 417 676 421
rect 682 421 686 425
rect 747 420 751 424
rect 757 420 761 424
rect 767 420 771 424
rect 777 424 781 428
rect 833 421 837 425
rect 843 442 847 446
rect 843 435 847 439
rect 859 421 863 425
rect 869 428 873 432
rect 879 436 883 440
rect 917 421 921 425
rect 927 442 931 446
rect 927 435 931 439
rect 943 421 947 425
rect 953 428 957 432
rect 1667 448 1671 452
rect 1717 461 1721 465
rect 1721 451 1725 455
rect 963 436 967 440
rect 979 420 983 424
rect 989 420 993 424
rect 999 420 1003 424
rect 1009 424 1013 428
rect 1721 441 1725 445
rect 1651 432 1655 436
rect 1721 431 1725 435
rect 1651 422 1655 426
rect 1651 412 1655 416
rect 1167 403 1171 407
rect 1200 403 1204 407
rect 1213 403 1217 407
rect 1230 403 1234 407
rect 1247 403 1251 407
rect 1267 403 1271 407
rect 1284 403 1288 407
rect 1301 403 1305 407
rect 1323 403 1327 407
rect 1340 403 1344 407
rect 1357 403 1361 407
rect 1377 403 1381 407
rect 1394 403 1398 407
rect 1411 403 1415 407
rect 1655 402 1659 406
rect 2034 398 2038 402
rect 2044 405 2048 409
rect 2044 398 2048 402
rect 2054 400 2058 404
rect 2064 412 2068 416
rect 2064 405 2068 409
rect 2121 398 2125 402
rect 2131 405 2135 409
rect 2131 398 2135 402
rect 2141 400 2145 404
rect 2151 412 2155 416
rect 2151 405 2155 409
rect 2214 398 2218 402
rect 2224 405 2228 409
rect 2224 398 2228 402
rect 2234 400 2238 404
rect 2244 412 2248 416
rect 2244 405 2248 409
rect 2454 414 2458 418
rect 2454 407 2458 411
rect 2547 414 2551 418
rect 2464 402 2468 406
rect 2474 407 2478 411
rect 2474 400 2478 404
rect 2547 407 2551 411
rect 2484 400 2488 404
rect 2634 414 2638 418
rect 2557 402 2561 406
rect 2567 407 2571 411
rect 2567 400 2571 404
rect 2634 407 2638 411
rect 2577 400 2581 404
rect 2644 402 2648 406
rect 2654 407 2658 411
rect 2654 400 2658 404
rect 2664 400 2668 404
rect 184 320 188 324
rect 1078 357 1082 361
rect 1122 357 1128 363
rect 1161 357 1165 361
rect 1194 357 1198 361
rect 1207 357 1211 361
rect 1224 357 1228 361
rect 1241 357 1245 361
rect 1261 357 1265 361
rect 1278 357 1282 361
rect 1295 357 1299 361
rect 1317 357 1321 361
rect 1334 357 1338 361
rect 1351 357 1355 361
rect 1371 357 1375 361
rect 1388 357 1392 361
rect 1405 357 1409 361
rect 214 322 218 326
rect 513 322 517 326
rect 202 313 206 317
rect 543 324 547 328
rect 840 325 844 329
rect 531 315 535 319
rect 870 327 874 331
rect 858 318 862 322
rect 1956 344 1960 348
rect 1966 344 1970 348
rect 1976 344 1980 348
rect 1986 348 1990 352
rect 1709 337 1713 341
rect 1713 327 1717 331
rect 90 269 94 273
rect 100 269 104 273
rect 110 269 114 273
rect 120 273 124 277
rect 176 270 180 274
rect 186 291 190 295
rect 186 284 190 288
rect 202 270 206 274
rect 212 277 216 281
rect 222 285 226 289
rect 260 270 264 274
rect 270 291 274 295
rect 270 284 274 288
rect 286 270 290 274
rect 296 277 300 281
rect 306 285 310 289
rect 322 269 326 273
rect 332 269 336 273
rect 342 269 346 273
rect 352 273 356 277
rect 419 271 423 275
rect 429 271 433 275
rect 439 271 443 275
rect 449 275 453 279
rect 505 272 509 276
rect 515 293 519 297
rect 515 286 519 290
rect 531 272 535 276
rect 541 279 545 283
rect 551 287 555 291
rect 589 272 593 276
rect 599 293 603 297
rect 599 286 603 290
rect 615 272 619 276
rect 625 279 629 283
rect 635 287 639 291
rect 651 271 655 275
rect 661 271 665 275
rect 671 271 675 275
rect 681 275 685 279
rect 746 274 750 278
rect 756 274 760 278
rect 766 274 770 278
rect 776 278 780 282
rect 832 275 836 279
rect 842 296 846 300
rect 842 289 846 293
rect 858 275 862 279
rect 868 282 872 286
rect 878 290 882 294
rect 916 275 920 279
rect 926 296 930 300
rect 926 289 930 293
rect 942 275 946 279
rect 952 282 956 286
rect 1452 302 1456 306
rect 962 290 966 294
rect 978 274 982 278
rect 988 274 992 278
rect 998 274 1002 278
rect 1008 278 1012 282
rect 1463 284 1467 288
rect 1713 317 1717 321
rect 2042 345 2046 349
rect 2052 366 2056 370
rect 2052 359 2056 363
rect 2068 345 2072 349
rect 2078 352 2082 356
rect 2088 360 2092 364
rect 2126 345 2130 349
rect 2136 366 2140 370
rect 2136 359 2140 363
rect 2152 345 2156 349
rect 2162 352 2166 356
rect 2172 360 2176 364
rect 2188 344 2192 348
rect 2198 344 2202 348
rect 2208 344 2212 348
rect 2218 348 2222 352
rect 2285 346 2289 350
rect 2295 346 2299 350
rect 2305 346 2309 350
rect 2315 350 2319 354
rect 1713 307 1717 311
rect 2371 347 2375 351
rect 2381 368 2385 372
rect 2381 361 2385 365
rect 2397 347 2401 351
rect 2407 354 2411 358
rect 2417 362 2421 366
rect 2455 347 2459 351
rect 2465 368 2469 372
rect 2465 361 2469 365
rect 2481 347 2485 351
rect 2491 354 2495 358
rect 2501 362 2505 366
rect 2517 346 2521 350
rect 2527 346 2531 350
rect 2537 346 2541 350
rect 2547 350 2551 354
rect 2612 349 2616 353
rect 2622 349 2626 353
rect 2632 349 2636 353
rect 2642 353 2646 357
rect 2698 350 2702 354
rect 2708 371 2712 375
rect 2708 364 2712 368
rect 2724 350 2728 354
rect 2734 357 2738 361
rect 2744 365 2748 369
rect 2782 350 2786 354
rect 2792 371 2796 375
rect 2792 364 2796 368
rect 2808 350 2812 354
rect 2818 357 2822 361
rect 2828 365 2832 369
rect 2844 349 2848 353
rect 2854 349 2858 353
rect 2864 349 2868 353
rect 2874 353 2878 357
rect 1474 301 1478 305
rect 1474 294 1478 298
rect 1697 291 1701 295
rect 1705 281 1709 285
rect 1712 271 1716 275
rect 1165 258 1169 262
rect 1198 258 1202 262
rect 1211 258 1215 262
rect 1228 258 1232 262
rect 1245 258 1249 262
rect 1265 258 1269 262
rect 1282 258 1286 262
rect 1299 258 1303 262
rect 1321 258 1325 262
rect 1338 258 1342 262
rect 1355 258 1359 262
rect 1375 258 1379 262
rect 1392 258 1396 262
rect 1409 258 1413 262
rect 1465 251 1469 255
rect 1691 255 1695 259
rect 1698 255 1702 259
rect 1454 233 1458 237
rect 183 174 187 178
rect 1079 215 1083 219
rect 1123 215 1129 221
rect 1476 241 1480 245
rect 1712 245 1716 249
rect 2049 249 2053 253
rect 1476 234 1480 238
rect 2079 251 2083 255
rect 2378 251 2382 255
rect 2067 242 2071 246
rect 2408 253 2412 257
rect 2705 254 2709 258
rect 2396 244 2400 248
rect 2735 256 2739 260
rect 2723 247 2727 251
rect 1162 215 1166 219
rect 1195 215 1199 219
rect 1208 215 1212 219
rect 1225 215 1229 219
rect 1242 215 1246 219
rect 1262 215 1266 219
rect 1279 215 1283 219
rect 1296 215 1300 219
rect 1318 215 1322 219
rect 1335 215 1339 219
rect 1352 215 1356 219
rect 1372 215 1376 219
rect 1389 215 1393 219
rect 1406 215 1410 219
rect 213 176 217 180
rect 512 176 516 180
rect 201 167 205 171
rect 542 178 546 182
rect 839 179 843 183
rect 530 169 534 173
rect 869 181 873 185
rect 1697 207 1701 211
rect 857 172 861 176
rect 1705 197 1709 201
rect 1712 187 1716 191
rect 1691 171 1695 175
rect 1698 171 1702 175
rect 384 129 388 133
rect 384 122 388 126
rect 394 134 398 138
rect 404 136 408 140
rect 404 129 408 133
rect 414 136 418 140
rect 477 129 481 133
rect 477 122 481 126
rect 487 134 491 138
rect 497 136 501 140
rect 497 129 501 133
rect 507 136 511 140
rect 564 129 568 133
rect 564 122 568 126
rect 574 134 578 138
rect 584 136 588 140
rect 584 129 588 133
rect 594 136 598 140
rect 1712 161 1716 165
rect 1806 198 1810 202
rect 1955 198 1959 202
rect 1965 198 1969 202
rect 1975 198 1979 202
rect 1985 202 1989 206
rect 1815 186 1819 190
rect 2041 199 2045 203
rect 2051 220 2055 224
rect 2051 213 2055 217
rect 2067 199 2071 203
rect 2077 206 2081 210
rect 2087 214 2091 218
rect 2125 199 2129 203
rect 2135 220 2139 224
rect 2135 213 2139 217
rect 2151 199 2155 203
rect 2161 206 2165 210
rect 2171 214 2175 218
rect 2187 198 2191 202
rect 2197 198 2201 202
rect 2207 198 2211 202
rect 2217 202 2221 206
rect 2284 200 2288 204
rect 2294 200 2298 204
rect 2304 200 2308 204
rect 2314 204 2318 208
rect 1808 168 1812 172
rect 2370 201 2374 205
rect 2380 222 2384 226
rect 2380 215 2384 219
rect 2396 201 2400 205
rect 2406 208 2410 212
rect 2416 216 2420 220
rect 2454 201 2458 205
rect 2464 222 2468 226
rect 2464 215 2468 219
rect 2480 201 2484 205
rect 2490 208 2494 212
rect 2500 216 2504 220
rect 2516 200 2520 204
rect 2526 200 2530 204
rect 2536 200 2540 204
rect 2546 204 2550 208
rect 2611 203 2615 207
rect 2621 203 2625 207
rect 2631 203 2635 207
rect 2641 207 2645 211
rect 2697 204 2701 208
rect 2707 225 2711 229
rect 2707 218 2711 222
rect 2723 204 2727 208
rect 2733 211 2737 215
rect 2743 219 2747 223
rect 2781 204 2785 208
rect 2791 225 2795 229
rect 2791 218 2795 222
rect 2807 204 2811 208
rect 2817 211 2821 215
rect 2827 219 2831 223
rect 2843 203 2847 207
rect 2853 203 2857 207
rect 2863 203 2867 207
rect 2873 207 2877 211
rect 1795 150 1799 154
rect 1802 150 1806 154
rect 1456 123 1460 127
rect 1166 116 1170 120
rect 1199 116 1203 120
rect 1212 116 1216 120
rect 1229 116 1233 120
rect 1246 116 1250 120
rect 1266 116 1270 120
rect 1283 116 1287 120
rect 1300 116 1304 120
rect 1322 116 1326 120
rect 1339 116 1343 120
rect 1356 116 1360 120
rect 1376 116 1380 120
rect 1393 116 1397 120
rect 1410 116 1414 120
rect 1467 105 1471 109
rect 1815 139 1819 143
rect 1478 122 1482 126
rect 1478 115 1482 119
rect 1795 127 1799 131
rect 1709 105 1713 109
rect 1713 95 1717 99
rect 1807 104 1811 108
rect 1814 104 1818 108
rect 2048 103 2052 107
rect 1799 92 1803 96
rect 1806 92 1810 96
rect 2078 105 2082 109
rect 2377 105 2381 109
rect 2066 96 2070 100
rect 2407 107 2411 111
rect 2704 108 2708 112
rect 2395 98 2399 102
rect 2734 110 2738 114
rect 2722 101 2726 105
rect 1713 85 1717 89
rect 1807 82 1811 86
rect 1814 82 1818 86
rect 1713 75 1717 79
rect 1792 72 1796 76
rect 1799 72 1803 76
rect 2249 58 2253 62
rect 2249 51 2253 55
rect 2259 63 2263 67
rect 2269 65 2273 69
rect 2269 58 2273 62
rect 2279 65 2283 69
rect 2342 58 2346 62
rect 2342 51 2346 55
rect 2352 63 2356 67
rect 2362 65 2366 69
rect 2362 58 2366 62
rect 2372 65 2376 69
rect 2429 58 2433 62
rect 2429 51 2433 55
rect 2439 63 2443 67
rect 2449 65 2453 69
rect 2449 58 2453 62
rect 2459 65 2463 69
<< m2contact >>
rect 1549 1101 1555 1107
rect 1813 1105 1817 1110
rect 1912 1105 1916 1111
rect 1921 1097 1925 1101
rect 1600 1072 1605 1080
rect 517 1041 522 1047
rect 153 1032 158 1037
rect 506 1035 510 1039
rect 989 1034 994 1039
rect 1042 1025 1046 1029
rect 505 1020 510 1025
rect 541 1020 546 1025
rect 75 1014 80 1020
rect 153 1008 157 1012
rect 145 982 150 987
rect 241 1008 245 1012
rect 237 982 241 986
rect 334 1008 338 1012
rect 382 1013 386 1017
rect 558 1013 563 1018
rect 286 981 290 985
rect 330 982 334 986
rect 1023 1021 1027 1025
rect 455 1001 460 1006
rect 516 1002 521 1007
rect 612 1010 616 1014
rect 382 990 386 994
rect 559 990 564 995
rect 616 984 620 988
rect 382 973 386 977
rect 560 973 564 977
rect 647 983 651 988
rect 705 1009 709 1013
rect 1068 1025 1072 1029
rect 792 1009 796 1013
rect 709 984 713 988
rect 722 986 726 990
rect 275 956 279 960
rect 312 957 317 961
rect 623 962 628 967
rect 658 962 662 967
rect 721 962 725 966
rect 735 961 739 965
rect 745 986 749 990
rect 987 992 993 998
rect 1090 998 1094 1002
rect 1162 997 1166 1001
rect 797 984 802 988
rect 745 962 749 966
rect 1105 988 1109 992
rect 1165 987 1169 991
rect 1187 997 1191 1001
rect 1209 998 1213 1002
rect 1177 987 1181 991
rect 1229 1005 1233 1009
rect 1239 997 1243 1001
rect 1206 983 1210 987
rect 1263 988 1267 992
rect 1296 997 1300 1001
rect 1332 1000 1336 1004
rect 1295 989 1299 993
rect 1312 992 1316 996
rect 1322 990 1326 994
rect 1285 982 1289 986
rect 1371 998 1375 1002
rect 1385 991 1389 995
rect 1354 983 1358 987
rect 103 936 107 940
rect 246 936 250 940
rect 79 908 83 912
rect 111 910 115 914
rect 148 910 152 914
rect 168 909 172 913
rect 304 927 308 931
rect 215 909 219 913
rect 252 909 256 913
rect 335 936 339 940
rect 350 927 354 931
rect 365 927 369 931
rect 304 893 308 897
rect 343 911 347 915
rect 60 882 64 886
rect 345 883 351 889
rect 172 841 176 845
rect 163 833 167 837
rect 365 859 369 863
rect 432 938 436 942
rect 461 929 465 934
rect 408 910 412 914
rect 440 912 444 916
rect 453 898 457 903
rect 575 938 579 942
rect 477 912 481 916
rect 497 911 501 915
rect 632 931 636 935
rect 544 911 548 915
rect 581 911 585 915
rect 664 938 668 942
rect 633 895 637 899
rect 672 913 676 917
rect 385 882 392 889
rect 672 885 678 891
rect 622 871 627 876
rect 390 859 394 863
rect 462 859 466 863
rect 501 843 505 847
rect 492 835 496 839
rect 684 856 688 860
rect 345 811 350 815
rect 365 810 370 815
rect 102 790 106 794
rect 759 941 763 945
rect 902 941 906 945
rect 794 931 798 935
rect 735 913 739 917
rect 767 915 771 919
rect 804 915 808 919
rect 824 914 828 918
rect 879 933 883 937
rect 871 914 875 918
rect 795 898 799 902
rect 880 898 884 902
rect 957 934 962 938
rect 908 914 912 918
rect 991 941 995 945
rect 960 898 964 902
rect 999 916 1003 920
rect 1181 940 1185 944
rect 1129 934 1134 939
rect 712 884 719 891
rect 796 868 801 873
rect 716 856 720 860
rect 787 856 791 860
rect 809 861 813 865
rect 828 846 832 850
rect 819 838 823 842
rect 872 861 876 865
rect 880 855 884 860
rect 809 830 813 834
rect 797 824 801 828
rect 879 820 884 827
rect 1166 930 1170 934
rect 1267 939 1271 943
rect 1299 938 1303 942
rect 1191 930 1195 934
rect 1213 930 1217 934
rect 1243 930 1247 934
rect 1326 937 1330 941
rect 1300 930 1304 934
rect 1358 944 1362 948
rect 1389 936 1393 940
rect 1336 927 1340 931
rect 1375 929 1379 933
rect 1233 922 1237 926
rect 1127 901 1132 906
rect 1729 1054 1733 1058
rect 1602 1047 1606 1051
rect 1704 1046 1708 1050
rect 1636 1025 1640 1029
rect 1603 951 1607 955
rect 1664 1001 1668 1005
rect 1719 1013 1723 1017
rect 1747 1015 1751 1019
rect 1638 993 1642 997
rect 1623 979 1628 984
rect 1664 979 1668 983
rect 1638 956 1642 960
rect 1561 941 1565 945
rect 1569 932 1573 936
rect 1637 936 1641 940
rect 1808 982 1812 986
rect 1731 963 1735 967
rect 1704 957 1708 961
rect 1703 937 1707 941
rect 1746 938 1750 942
rect 1151 883 1155 887
rect 1090 853 1094 857
rect 1162 852 1166 856
rect 1105 843 1109 847
rect 1187 852 1191 856
rect 1209 852 1213 856
rect 1229 860 1233 864
rect 1239 852 1243 856
rect 1177 842 1181 846
rect 1263 843 1267 847
rect 1296 852 1300 856
rect 1332 855 1336 859
rect 1295 844 1299 848
rect 1312 847 1316 851
rect 1322 845 1326 849
rect 1285 837 1289 841
rect 1371 853 1375 857
rect 1385 846 1389 850
rect 1354 838 1358 842
rect 998 820 1002 824
rect 78 762 82 766
rect 110 764 114 768
rect 147 764 151 768
rect 167 763 171 767
rect 214 763 218 767
rect 245 790 249 794
rect 334 790 338 794
rect 351 782 355 786
rect 251 763 255 767
rect 303 771 307 775
rect 228 747 232 751
rect 303 747 307 751
rect 342 765 346 769
rect 345 737 353 744
rect 294 727 298 731
rect 364 728 368 732
rect 171 695 175 699
rect 162 687 166 691
rect 289 708 295 714
rect 318 708 323 713
rect 343 708 348 713
rect 364 708 369 713
rect 431 792 435 796
rect 574 792 578 796
rect 467 773 471 777
rect 407 764 411 768
rect 439 766 443 770
rect 476 766 480 770
rect 496 765 500 769
rect 543 765 547 769
rect 467 749 471 753
rect 632 777 636 781
rect 663 792 667 796
rect 580 765 584 769
rect 632 749 636 753
rect 671 767 675 771
rect 382 737 387 742
rect 672 738 676 742
rect 391 728 395 732
rect 467 723 471 727
rect 467 705 471 709
rect 426 675 430 679
rect 500 697 504 701
rect 491 689 495 693
rect 557 715 563 720
rect 645 715 650 720
rect 540 682 545 687
rect 439 675 443 679
rect 428 661 432 665
rect 450 661 454 665
rect 628 660 632 665
rect 439 646 443 650
rect 411 609 416 614
rect 431 598 435 602
rect 541 638 545 643
rect 508 626 512 631
rect 504 609 509 614
rect 597 626 601 630
rect 758 795 762 799
rect 901 795 905 799
rect 734 767 738 771
rect 766 769 770 773
rect 803 769 807 773
rect 823 768 827 772
rect 870 768 874 772
rect 959 779 963 783
rect 990 795 994 799
rect 907 768 911 772
rect 959 752 963 756
rect 998 770 1002 774
rect 712 738 716 742
rect 770 729 774 733
rect 709 715 714 720
rect 743 715 748 720
rect 827 700 831 704
rect 818 692 822 696
rect 875 717 881 722
rect 770 688 774 692
rect 1391 822 1395 826
rect 1181 795 1185 799
rect 1166 785 1170 789
rect 1267 794 1271 798
rect 1299 793 1303 797
rect 1191 785 1195 789
rect 1213 785 1217 789
rect 1243 785 1247 789
rect 1326 792 1330 796
rect 1300 785 1304 789
rect 1358 799 1362 803
rect 1389 791 1393 795
rect 1336 782 1340 786
rect 1375 784 1379 788
rect 1233 777 1237 781
rect 1462 886 1469 892
rect 1413 861 1417 865
rect 1562 891 1566 895
rect 1557 874 1564 880
rect 1637 889 1641 893
rect 1731 926 1735 930
rect 1768 937 1772 941
rect 1412 823 1416 827
rect 1469 819 1474 825
rect 1415 782 1419 786
rect 1447 783 1451 787
rect 1093 742 1097 746
rect 1148 738 1152 742
rect 1089 711 1093 715
rect 1161 710 1165 714
rect 1104 701 1108 705
rect 1186 710 1190 714
rect 1208 710 1212 714
rect 1228 718 1232 722
rect 1238 710 1242 714
rect 1176 700 1180 704
rect 1262 701 1266 705
rect 1295 710 1299 714
rect 1331 713 1335 717
rect 1294 702 1298 706
rect 1311 705 1315 709
rect 1321 703 1325 707
rect 1284 695 1288 699
rect 1370 711 1374 715
rect 1384 704 1388 708
rect 1353 696 1357 700
rect 720 653 725 659
rect 1050 632 1054 636
rect 1052 622 1058 628
rect 1033 618 1037 622
rect 589 609 594 614
rect 1042 610 1046 614
rect 1180 653 1184 657
rect 1165 643 1169 647
rect 1102 629 1106 633
rect 1266 652 1270 656
rect 1298 651 1302 655
rect 1190 643 1194 647
rect 1212 643 1216 647
rect 1242 643 1246 647
rect 1325 650 1329 654
rect 1299 643 1303 647
rect 1357 657 1361 661
rect 1388 649 1392 653
rect 1335 640 1339 644
rect 1374 642 1378 646
rect 1232 635 1236 639
rect 1101 614 1105 618
rect 1134 613 1139 617
rect 1396 613 1400 617
rect 1415 711 1419 715
rect 1446 716 1450 720
rect 1438 675 1443 679
rect 1664 858 1668 862
rect 1637 852 1641 856
rect 1594 823 1599 828
rect 1583 813 1588 818
rect 1553 787 1558 792
rect 1554 773 1559 778
rect 1602 810 1606 814
rect 1602 788 1606 792
rect 1731 879 1735 883
rect 1799 883 1803 887
rect 1807 874 1811 878
rect 1730 859 1734 863
rect 1730 822 1734 826
rect 1621 800 1625 804
rect 1647 800 1651 804
rect 1704 814 1708 818
rect 1787 838 1791 842
rect 1815 836 1820 840
rect 1732 790 1736 794
rect 1664 769 1668 773
rect 1760 767 1768 775
rect 1639 761 1643 765
rect 1553 727 1558 732
rect 1768 741 1772 745
rect 1733 722 1740 728
rect 1564 711 1569 716
rect 1590 712 1595 717
rect 1422 603 1427 607
rect 225 584 230 591
rect 355 587 362 594
rect 1091 589 1096 594
rect 1458 603 1462 607
rect 1019 558 1026 563
rect 1041 558 1047 564
rect 528 535 533 541
rect 164 526 169 531
rect 86 508 91 514
rect 164 502 168 506
rect 156 476 161 481
rect 252 502 256 506
rect 248 476 252 480
rect 345 502 349 506
rect 393 507 397 511
rect 466 507 472 513
rect 569 507 574 512
rect 297 475 301 479
rect 341 476 345 480
rect 474 497 478 502
rect 527 496 532 501
rect 393 484 397 488
rect 454 485 460 491
rect 623 504 627 508
rect 570 485 575 489
rect 435 474 441 480
rect 529 475 534 480
rect 556 475 561 480
rect 627 478 631 482
rect 393 467 397 471
rect 571 467 575 471
rect 658 477 662 482
rect 716 503 720 507
rect 803 503 807 507
rect 1062 573 1066 577
rect 1096 566 1100 570
rect 1152 568 1157 573
rect 1057 558 1064 566
rect 1174 557 1182 564
rect 1142 546 1147 550
rect 1150 512 1155 517
rect 720 478 724 482
rect 733 480 737 484
rect 286 450 290 454
rect 323 451 328 455
rect 634 456 639 461
rect 669 456 673 461
rect 732 456 736 460
rect 746 455 750 459
rect 756 480 760 484
rect 808 478 813 482
rect 756 456 760 460
rect 1033 489 1037 494
rect 1082 489 1087 493
rect 1111 487 1115 491
rect 1183 486 1187 490
rect 1126 477 1130 481
rect 1208 486 1212 490
rect 1230 486 1234 490
rect 1250 494 1254 498
rect 1260 486 1264 490
rect 1198 476 1202 480
rect 1284 477 1288 481
rect 1317 486 1321 490
rect 1353 489 1357 493
rect 1316 478 1320 482
rect 1333 481 1337 485
rect 1343 479 1347 483
rect 1306 471 1310 475
rect 1392 487 1396 491
rect 1406 480 1410 484
rect 1375 472 1379 476
rect 114 430 118 434
rect 257 430 261 434
rect 90 402 94 406
rect 122 404 126 408
rect 159 404 163 408
rect 179 403 183 407
rect 226 403 230 407
rect 346 431 350 435
rect 360 422 364 426
rect 263 403 267 407
rect 315 411 319 415
rect 315 387 319 391
rect 354 405 358 409
rect 71 376 75 380
rect 356 377 362 383
rect 345 363 350 368
rect 183 335 187 339
rect 174 327 178 331
rect 376 353 380 357
rect 443 432 447 436
rect 586 432 590 436
rect 419 404 423 408
rect 451 406 455 410
rect 488 406 492 410
rect 508 405 512 409
rect 643 425 647 429
rect 555 405 559 409
rect 592 405 596 409
rect 675 432 679 436
rect 644 389 648 393
rect 683 407 687 411
rect 396 376 403 383
rect 683 379 689 385
rect 487 365 492 370
rect 401 353 405 357
rect 473 353 477 357
rect 344 325 349 331
rect 376 325 380 330
rect 583 365 588 370
rect 672 365 677 369
rect 512 337 516 341
rect 486 325 491 330
rect 503 329 507 333
rect 695 350 699 354
rect 672 333 676 337
rect 770 435 774 439
rect 913 435 917 439
rect 805 425 809 429
rect 790 417 794 421
rect 746 407 750 411
rect 778 409 782 413
rect 788 393 792 398
rect 815 409 819 413
rect 835 408 839 412
rect 890 427 894 431
rect 882 408 886 412
rect 806 392 810 396
rect 891 392 895 396
rect 968 428 973 432
rect 919 408 923 412
rect 1002 435 1006 439
rect 971 392 975 396
rect 1010 410 1014 414
rect 723 378 730 385
rect 356 305 361 309
rect 376 304 381 309
rect 113 284 117 288
rect 89 256 93 260
rect 121 258 125 262
rect 158 258 162 262
rect 178 257 182 261
rect 225 257 229 261
rect 256 284 260 288
rect 314 272 318 276
rect 262 257 266 261
rect 239 241 243 245
rect 345 284 349 288
rect 361 276 365 280
rect 376 276 380 280
rect 314 241 318 245
rect 353 259 357 263
rect 356 231 364 238
rect 305 221 309 225
rect 182 189 186 193
rect 173 181 177 185
rect 300 202 306 208
rect 329 202 334 207
rect 336 178 340 182
rect 354 202 359 207
rect 375 202 380 207
rect 442 286 446 290
rect 585 286 589 290
rect 478 267 482 271
rect 418 258 422 262
rect 450 260 454 264
rect 487 260 491 264
rect 507 259 511 263
rect 554 259 558 263
rect 478 243 482 247
rect 643 270 647 274
rect 674 286 678 290
rect 591 259 595 263
rect 643 243 647 247
rect 682 261 686 265
rect 393 231 398 236
rect 683 232 687 236
rect 427 223 431 228
rect 489 225 493 229
rect 478 217 482 221
rect 402 210 406 215
rect 454 210 458 215
rect 427 201 432 207
rect 631 225 635 229
rect 355 178 360 183
rect 375 178 380 183
rect 428 168 432 173
rect 478 199 482 203
rect 511 191 515 195
rect 502 183 506 187
rect 568 209 574 214
rect 656 209 661 214
rect 675 190 680 194
rect 551 176 556 181
rect 450 169 454 173
rect 755 359 760 364
rect 807 362 812 367
rect 727 350 731 354
rect 798 350 802 354
rect 820 355 824 359
rect 839 340 843 344
rect 830 332 834 336
rect 883 355 887 359
rect 891 349 895 354
rect 1062 437 1068 443
rect 1202 429 1206 433
rect 1187 419 1191 423
rect 1288 428 1292 432
rect 1320 427 1324 431
rect 1212 419 1216 423
rect 1234 419 1238 423
rect 1264 419 1268 423
rect 1347 426 1351 430
rect 1321 419 1325 423
rect 1379 433 1383 437
rect 1410 425 1414 429
rect 1357 416 1361 420
rect 1396 418 1400 422
rect 1254 411 1258 415
rect 1062 392 1068 398
rect 1449 437 1455 443
rect 1171 372 1175 376
rect 820 324 824 328
rect 739 317 743 322
rect 808 318 812 322
rect 890 314 895 321
rect 1003 312 1007 317
rect 1109 342 1113 346
rect 1181 341 1185 345
rect 1124 332 1128 336
rect 1206 341 1210 345
rect 1228 341 1232 345
rect 1248 349 1252 353
rect 1258 341 1262 345
rect 1196 331 1200 335
rect 1282 332 1286 336
rect 1315 341 1319 345
rect 1351 344 1355 348
rect 1314 333 1318 337
rect 1331 336 1335 340
rect 1341 334 1345 338
rect 1304 326 1308 330
rect 1390 342 1394 346
rect 1404 335 1408 339
rect 1373 327 1377 331
rect 769 289 773 293
rect 794 280 798 285
rect 745 261 749 265
rect 777 263 781 267
rect 912 289 916 293
rect 814 263 818 267
rect 834 262 838 266
rect 881 262 885 266
rect 792 250 796 255
rect 970 273 974 277
rect 1001 289 1005 293
rect 918 262 922 266
rect 970 246 974 250
rect 1009 264 1013 268
rect 723 232 727 236
rect 781 223 785 227
rect 720 209 725 214
rect 754 209 759 214
rect 781 182 785 186
rect 797 201 801 205
rect 886 211 892 216
rect 838 194 842 198
rect 829 186 833 190
rect 796 177 800 182
rect 1411 305 1415 309
rect 1365 298 1369 302
rect 1200 284 1204 288
rect 1185 274 1189 278
rect 1286 283 1290 287
rect 1318 282 1322 286
rect 1210 274 1214 278
rect 1232 274 1236 278
rect 1262 274 1266 278
rect 1345 281 1349 285
rect 1319 274 1323 278
rect 1355 271 1359 275
rect 1252 266 1256 270
rect 1377 288 1381 292
rect 1408 280 1412 284
rect 1394 273 1398 277
rect 1564 682 1568 686
rect 1580 685 1584 689
rect 1580 659 1584 663
rect 1731 694 1735 698
rect 1706 686 1710 690
rect 1767 701 1772 705
rect 1638 665 1642 669
rect 1595 644 1599 648
rect 1666 641 1670 645
rect 1721 655 1725 659
rect 1749 655 1753 659
rect 1640 633 1644 637
rect 1623 622 1628 627
rect 1649 622 1654 627
rect 1627 612 1631 616
rect 1648 608 1652 612
rect 1640 596 1644 600
rect 1563 581 1567 585
rect 1571 572 1575 576
rect 1639 576 1643 580
rect 1733 603 1737 607
rect 1706 597 1710 601
rect 1705 577 1709 581
rect 1748 578 1752 582
rect 1580 540 1584 544
rect 1639 529 1643 533
rect 1733 566 1737 570
rect 1770 577 1774 581
rect 1624 516 1628 520
rect 1648 516 1652 520
rect 1666 498 1670 502
rect 1639 492 1643 496
rect 1489 468 1495 474
rect 1490 438 1496 444
rect 1531 437 1537 443
rect 1444 314 1448 318
rect 1489 309 1493 315
rect 1435 294 1439 298
rect 1365 245 1369 249
rect 1170 229 1174 233
rect 1110 200 1114 204
rect 1182 199 1186 203
rect 1125 190 1129 194
rect 1207 199 1211 203
rect 1229 199 1233 203
rect 1249 207 1253 211
rect 1259 199 1263 203
rect 1197 189 1201 193
rect 1283 190 1287 194
rect 1364 214 1368 218
rect 1316 199 1320 203
rect 1352 202 1356 206
rect 1315 191 1319 195
rect 1332 194 1336 198
rect 1342 192 1346 196
rect 1305 184 1309 188
rect 1391 200 1395 204
rect 1405 193 1409 197
rect 1374 185 1378 189
rect 1361 175 1365 179
rect 766 152 771 158
rect 450 140 454 144
rect 374 104 379 109
rect 422 103 427 108
rect 442 92 446 96
rect 552 132 556 137
rect 519 120 523 125
rect 515 103 520 108
rect 1052 128 1056 132
rect 608 120 612 124
rect 600 103 605 108
rect 366 81 373 88
rect 1412 163 1416 167
rect 1110 153 1114 157
rect 1148 153 1152 158
rect 1364 156 1368 160
rect 1201 142 1205 146
rect 1186 132 1190 136
rect 1287 141 1291 145
rect 1319 140 1323 144
rect 1211 132 1215 136
rect 1233 132 1237 136
rect 1263 132 1267 136
rect 1346 139 1350 143
rect 1320 132 1324 136
rect 1356 129 1360 133
rect 1253 124 1257 128
rect 1378 146 1382 150
rect 1409 138 1413 142
rect 1395 131 1399 135
rect 1365 101 1369 105
rect 1447 224 1451 228
rect 1589 457 1593 461
rect 1560 348 1565 354
rect 1510 328 1514 332
rect 1600 450 1604 454
rect 1733 519 1737 523
rect 1801 523 1805 527
rect 1809 514 1813 518
rect 1732 499 1736 503
rect 1770 493 1778 502
rect 1732 462 1736 466
rect 1623 440 1627 444
rect 1649 440 1653 444
rect 1706 454 1710 458
rect 1782 479 1788 485
rect 1818 478 1824 484
rect 1734 430 1738 434
rect 1810 431 1816 437
rect 1666 409 1670 413
rect 1762 407 1770 415
rect 1641 401 1645 405
rect 1684 398 1690 404
rect 1709 384 1715 391
rect 1758 381 1765 389
rect 1808 382 1814 387
rect 1735 362 1742 368
rect 1685 350 1690 355
rect 1772 353 1776 357
rect 1801 353 1805 357
rect 1723 338 1727 342
rect 1600 320 1604 325
rect 1698 330 1702 334
rect 1506 292 1510 298
rect 1645 288 1650 294
rect 1770 317 1777 324
rect 1710 299 1714 303
rect 1741 299 1745 303
rect 1488 221 1492 225
rect 1504 221 1508 225
rect 1647 220 1651 224
rect 1447 170 1451 174
rect 1440 139 1444 143
rect 1488 135 1492 139
rect 1922 1082 1926 1087
rect 1903 989 1908 998
rect 1944 1097 1948 1103
rect 1929 963 1933 967
rect 2006 1082 2013 1087
rect 2005 924 2009 928
rect 2083 889 2087 894
rect 2631 982 2635 986
rect 2708 974 2712 978
rect 2799 966 2803 970
rect 2708 962 2712 966
rect 2800 945 2804 949
rect 2631 935 2635 939
rect 2288 924 2292 928
rect 2210 888 2214 892
rect 2451 892 2455 896
rect 2492 909 2496 913
rect 2877 924 2881 928
rect 2788 918 2792 922
rect 2483 901 2487 905
rect 2570 892 2574 896
rect 2596 892 2600 896
rect 2379 879 2384 883
rect 2380 869 2384 873
rect 1818 307 1822 311
rect 1780 289 1784 293
rect 1905 768 1911 776
rect 2005 848 2010 854
rect 2210 848 2214 852
rect 2131 819 2136 823
rect 2132 795 2136 799
rect 2211 795 2215 799
rect 1940 766 1944 772
rect 1963 776 1968 781
rect 1959 743 1966 747
rect 2009 774 2013 778
rect 2055 766 2059 770
rect 1985 746 1989 750
rect 2017 748 2021 752
rect 2054 748 2058 752
rect 2074 747 2078 751
rect 2121 747 2125 751
rect 2152 774 2156 778
rect 2210 782 2214 786
rect 2261 786 2266 791
rect 2241 774 2245 778
rect 2158 747 2162 751
rect 2131 731 2135 735
rect 2210 731 2214 735
rect 2249 749 2253 753
rect 2312 831 2316 835
rect 2351 849 2355 853
rect 2320 806 2324 810
rect 2354 824 2358 828
rect 2403 833 2407 837
rect 2440 833 2444 837
rect 2487 833 2491 837
rect 2507 832 2511 836
rect 2544 832 2548 836
rect 2576 834 2580 838
rect 2409 806 2413 810
rect 2552 806 2556 810
rect 2674 899 2678 903
rect 2718 894 2722 898
rect 2763 887 2767 891
rect 2807 910 2811 914
rect 2807 895 2811 899
rect 2852 911 2856 915
rect 2843 903 2847 907
rect 2877 894 2881 898
rect 2868 887 2872 891
rect 2951 887 2955 891
rect 2787 870 2791 874
rect 2850 878 2854 882
rect 2951 878 2955 882
rect 2309 786 2315 792
rect 2273 734 2279 741
rect 2295 761 2302 767
rect 1994 705 1998 709
rect 2078 679 2082 683
rect 2069 671 2073 675
rect 2225 680 2230 684
rect 2065 663 2069 667
rect 2292 711 2300 718
rect 2293 662 2298 668
rect 2365 766 2369 770
rect 2488 767 2492 771
rect 2401 750 2406 756
rect 2341 738 2345 742
rect 2373 740 2377 744
rect 2410 740 2414 744
rect 2401 732 2405 736
rect 2430 739 2434 743
rect 2477 739 2481 743
rect 2508 766 2512 770
rect 2566 749 2570 753
rect 2597 766 2601 770
rect 2514 739 2518 743
rect 2489 724 2493 728
rect 2566 723 2570 727
rect 2605 741 2609 745
rect 2672 833 2676 837
rect 2711 851 2715 855
rect 2780 851 2786 855
rect 2763 835 2767 839
rect 2680 808 2684 812
rect 2712 823 2716 827
rect 2800 835 2804 839
rect 2787 824 2791 828
rect 2847 835 2851 839
rect 2867 834 2871 838
rect 2904 834 2908 838
rect 2936 836 2940 840
rect 2769 808 2773 812
rect 2912 808 2916 812
rect 2633 736 2639 743
rect 2318 706 2326 714
rect 2488 702 2492 706
rect 2401 685 2406 690
rect 1902 633 1908 639
rect 1927 619 1935 624
rect 1911 606 1920 611
rect 1928 568 1934 574
rect 1902 516 1908 522
rect 1943 538 1952 546
rect 2268 641 2272 645
rect 2342 660 2348 666
rect 2434 671 2438 675
rect 2402 658 2407 664
rect 2425 663 2429 667
rect 2725 768 2729 772
rect 2848 769 2852 773
rect 2751 752 2755 756
rect 2701 740 2705 744
rect 2733 742 2737 746
rect 2770 742 2774 746
rect 2790 741 2794 745
rect 2837 741 2841 745
rect 2752 731 2756 735
rect 2762 731 2766 735
rect 2868 768 2872 772
rect 2874 741 2878 745
rect 2925 749 2929 754
rect 2957 768 2961 772
rect 2849 726 2853 730
rect 2926 725 2930 729
rect 2965 743 2969 747
rect 2678 708 2686 716
rect 2752 694 2757 700
rect 2848 704 2852 708
rect 2762 680 2767 686
rect 2754 662 2759 668
rect 2794 673 2798 677
rect 2763 661 2768 667
rect 2785 665 2789 669
rect 2019 636 2023 640
rect 2064 634 2068 638
rect 1994 628 1998 632
rect 2619 625 2623 629
rect 2034 585 2039 589
rect 2262 567 2266 571
rect 2245 490 2251 495
rect 1982 476 1986 481
rect 2197 477 2202 482
rect 2909 507 2913 511
rect 2393 464 2398 470
rect 1951 437 1956 443
rect 1981 458 1985 462
rect 1915 422 1920 428
rect 1897 414 1902 418
rect 1962 413 1967 419
rect 2029 455 2034 460
rect 2197 454 2202 461
rect 1995 432 1999 437
rect 2029 431 2033 435
rect 2021 405 2026 410
rect 2117 431 2121 435
rect 2113 405 2117 409
rect 2210 431 2214 435
rect 2258 436 2262 440
rect 2434 436 2439 441
rect 2162 404 2166 408
rect 2206 405 2210 409
rect 2293 427 2298 432
rect 2392 425 2397 430
rect 2488 433 2492 437
rect 2258 413 2262 417
rect 2435 413 2440 418
rect 2492 407 2496 411
rect 2258 396 2262 400
rect 2436 396 2440 400
rect 2523 406 2527 411
rect 2581 432 2585 436
rect 2668 432 2672 436
rect 2585 407 2589 411
rect 2598 409 2602 413
rect 2151 379 2155 383
rect 2188 380 2193 384
rect 2499 385 2504 390
rect 2534 385 2538 390
rect 2597 385 2601 389
rect 2611 384 2615 388
rect 2621 409 2625 413
rect 2673 407 2678 411
rect 2621 385 2625 389
rect 1725 247 1729 251
rect 1698 241 1702 245
rect 1741 220 1745 224
rect 1725 210 1729 214
rect 1768 246 1772 250
rect 1761 210 1765 214
rect 1874 274 1879 280
rect 1534 135 1538 139
rect 1498 106 1503 112
rect 1098 90 1103 95
rect 1581 91 1586 97
rect 1725 163 1729 167
rect 1777 167 1781 171
rect 1797 167 1801 171
rect 1724 143 1728 147
rect 1740 132 1744 136
rect 1764 159 1768 163
rect 1786 159 1790 163
rect 1724 106 1728 110
rect 1698 98 1702 102
rect 1808 141 1812 145
rect 1783 112 1787 116
rect 1626 79 1633 86
rect 1650 77 1655 82
rect 1674 77 1678 82
rect 1349 56 1356 62
rect 1650 56 1655 62
rect 983 44 992 53
rect 1528 43 1534 50
rect 1056 29 1063 37
rect 1621 26 1625 30
rect 1398 17 1403 22
rect 1516 18 1523 26
rect 1726 74 1730 78
rect 1767 83 1771 87
rect 1696 52 1701 57
rect 1735 52 1740 57
rect 1795 50 1799 55
rect 1697 30 1702 36
rect 1717 29 1723 34
rect 1736 32 1740 37
rect 1979 359 1983 363
rect 2122 359 2126 363
rect 1955 331 1959 335
rect 1987 333 1991 337
rect 2024 333 2028 337
rect 2044 332 2048 336
rect 2176 352 2180 356
rect 2091 332 2095 336
rect 2128 332 2132 336
rect 2211 359 2215 363
rect 2241 361 2245 366
rect 2180 316 2184 320
rect 2219 334 2223 338
rect 1936 305 1940 309
rect 2221 306 2227 312
rect 2242 294 2246 299
rect 2048 264 2052 268
rect 2039 256 2043 260
rect 2241 282 2245 286
rect 2308 361 2312 365
rect 2451 361 2455 365
rect 2284 333 2288 337
rect 2316 335 2320 339
rect 2353 335 2357 339
rect 2373 334 2377 338
rect 2508 354 2512 358
rect 2420 334 2424 338
rect 2457 334 2461 338
rect 2540 361 2544 365
rect 2509 318 2513 322
rect 2548 336 2552 340
rect 2261 305 2268 312
rect 2548 308 2554 314
rect 2259 294 2264 299
rect 2266 282 2270 286
rect 2338 282 2342 286
rect 2377 266 2381 270
rect 2267 258 2273 263
rect 2368 258 2372 262
rect 2560 279 2564 283
rect 2635 364 2639 368
rect 2778 364 2782 368
rect 2670 354 2674 358
rect 2611 336 2615 340
rect 2643 338 2647 342
rect 2680 338 2684 342
rect 2700 337 2704 341
rect 2755 356 2759 360
rect 2747 337 2751 341
rect 2671 321 2675 325
rect 2756 321 2760 325
rect 2833 357 2838 361
rect 2784 337 2788 341
rect 2867 364 2871 368
rect 2836 321 2840 325
rect 2875 339 2879 343
rect 2588 307 2595 314
rect 2672 291 2677 296
rect 2592 279 2596 283
rect 2663 279 2667 283
rect 2221 234 2226 238
rect 2241 233 2246 238
rect 2685 284 2689 288
rect 2704 269 2708 273
rect 2695 261 2699 265
rect 2748 284 2752 288
rect 2756 278 2760 283
rect 2685 253 2689 257
rect 2673 247 2677 251
rect 2755 243 2760 250
rect 2866 245 2870 249
rect 1978 213 1982 217
rect 1954 185 1958 189
rect 1986 187 1990 191
rect 2023 187 2027 191
rect 2043 186 2047 190
rect 2090 186 2094 190
rect 2121 213 2125 217
rect 2210 213 2214 217
rect 2127 186 2131 190
rect 2179 194 2183 198
rect 2104 170 2108 174
rect 2179 170 2183 174
rect 2218 188 2222 192
rect 2221 160 2229 167
rect 2170 150 2174 154
rect 2047 118 2051 122
rect 2038 110 2042 114
rect 2165 131 2171 137
rect 2194 131 2199 136
rect 1966 72 1970 77
rect 2219 131 2224 136
rect 2240 131 2245 136
rect 2307 215 2311 219
rect 2450 215 2454 219
rect 2343 196 2347 200
rect 2283 187 2287 191
rect 2315 189 2319 193
rect 2352 189 2356 193
rect 2372 188 2376 192
rect 2419 188 2423 192
rect 2343 172 2347 176
rect 2539 215 2543 219
rect 2456 188 2460 192
rect 2508 195 2512 199
rect 2508 172 2512 176
rect 2547 190 2551 194
rect 2258 160 2263 165
rect 2548 161 2552 165
rect 2343 146 2347 150
rect 2343 128 2347 132
rect 2376 120 2380 124
rect 2367 112 2371 116
rect 2433 138 2439 143
rect 2521 138 2526 143
rect 2634 218 2638 222
rect 2777 218 2781 222
rect 2835 226 2839 230
rect 2610 190 2614 194
rect 2642 192 2646 196
rect 2679 192 2683 196
rect 2699 191 2703 195
rect 2746 191 2750 195
rect 2866 218 2870 222
rect 2783 191 2787 195
rect 2835 198 2839 202
rect 2835 175 2839 179
rect 2874 193 2878 197
rect 2588 161 2592 165
rect 2646 152 2650 156
rect 2585 138 2590 143
rect 2619 138 2624 143
rect 2416 105 2421 110
rect 2315 98 2319 102
rect 2703 123 2707 127
rect 2694 115 2698 119
rect 2751 140 2757 145
rect 2646 111 2650 115
rect 2315 69 2319 73
rect 1772 26 1777 31
rect 1683 18 1688 23
rect 1706 8 1710 12
rect 1798 30 1802 34
rect 2287 32 2292 37
rect 1837 16 1843 22
rect 2307 21 2311 25
rect 2417 61 2421 66
rect 2384 49 2388 54
rect 2380 32 2385 37
rect 2473 49 2477 53
rect 2465 32 2470 37
rect 2231 10 2238 17
rect 1849 2 1856 10
rect 1878 -8 1884 -3
rect 2298 -8 2302 -4
<< m3contact >>
rect 541 958 545 962
rect 560 937 564 941
rect 326 589 332 596
rect 1478 887 1483 892
rect 1558 864 1563 869
rect 31 474 35 479
rect 568 476 572 480
rect 1202 709 1206 713
rect 1343 622 1348 627
rect 1057 612 1062 617
rect 552 452 556 456
rect 571 431 575 435
rect 699 395 703 400
rect 730 318 734 322
rect 459 211 464 217
rect 995 220 1000 224
rect 762 180 767 186
rect 730 176 734 180
rect 647 154 652 158
rect 952 170 958 176
rect 1344 567 1348 571
rect 1222 558 1228 565
rect 1225 486 1229 490
rect 1812 989 1817 994
rect 1820 953 1825 960
rect 1844 861 1850 869
rect 1223 341 1227 345
rect 1544 361 1550 367
rect 1786 495 1791 502
rect 1544 301 1549 307
rect 1084 248 1089 252
rect 1223 200 1227 204
rect 1640 278 1646 284
rect 1652 220 1657 226
rect 669 83 673 87
rect 954 46 959 52
rect 1581 44 1586 51
rect 1627 39 1633 45
rect 1645 26 1649 30
rect 1787 49 1791 53
rect 1761 27 1765 31
rect 1895 991 1899 995
rect 1886 955 1894 961
rect 1934 813 1942 822
rect 2023 640 2027 644
rect 2262 639 2266 643
rect 2023 585 2027 589
rect 2262 577 2266 581
rect 2182 538 2186 542
rect 2104 517 2108 521
rect 1904 435 1909 442
rect 2606 432 2610 436
rect 2180 400 2184 405
rect 2417 381 2421 385
rect 2103 353 2107 357
rect 2436 360 2440 364
rect 2007 244 2012 250
rect 1898 220 1902 224
rect 2179 200 2183 204
rect 2256 245 2261 251
rect 1941 73 1945 79
rect 1866 13 1873 19
rect 2507 203 2512 208
rect 1582 -10 1586 -3
<< psubstratepcontact >>
rect 187 1025 191 1029
rect 274 1025 278 1029
rect 367 1025 371 1029
rect 579 1027 583 1031
rect 672 1027 676 1031
rect 759 1027 763 1031
rect 1614 1023 1618 1027
rect 1754 1024 1758 1028
rect 81 886 85 890
rect 159 886 163 890
rect 243 886 247 890
rect 313 886 317 890
rect 410 888 414 892
rect 488 888 492 892
rect 572 888 576 892
rect 1754 954 1758 958
rect 1614 945 1618 949
rect 642 888 646 892
rect 737 891 741 895
rect 815 891 819 895
rect 899 891 903 895
rect 1604 930 1608 934
rect 1764 913 1768 917
rect 1604 902 1608 906
rect 969 891 973 895
rect 174 876 178 880
rect 202 876 206 880
rect 503 878 507 882
rect 531 878 535 882
rect 830 881 834 885
rect 858 881 862 885
rect 1764 885 1768 889
rect 1754 870 1758 874
rect 1614 861 1618 865
rect 2453 866 2457 870
rect 2481 866 2485 870
rect 2813 868 2817 872
rect 2841 868 2845 872
rect 2342 856 2346 860
rect 1421 826 1425 830
rect 2412 856 2416 860
rect 2496 856 2500 860
rect 2574 856 2578 860
rect 2702 858 2706 862
rect 1422 817 1426 821
rect 80 740 84 744
rect 158 740 162 744
rect 242 740 246 744
rect 312 740 316 744
rect 409 742 413 746
rect 487 742 491 746
rect 571 742 575 746
rect 1614 791 1618 795
rect 641 742 645 746
rect 736 745 740 749
rect 814 745 818 749
rect 898 745 902 749
rect 1754 792 1758 796
rect 2772 858 2776 862
rect 2856 858 2860 862
rect 2934 858 2938 862
rect 968 745 972 749
rect 173 730 177 734
rect 201 730 205 734
rect 502 732 506 736
rect 530 732 534 736
rect 829 735 833 739
rect 857 735 861 739
rect 1987 724 1991 728
rect 2065 724 2069 728
rect 2149 724 2153 728
rect 2219 724 2223 728
rect 1421 686 1425 690
rect 2080 714 2084 718
rect 2108 714 2112 718
rect 2343 716 2347 720
rect 2421 716 2425 720
rect 2505 716 2509 720
rect 2575 716 2579 720
rect 2703 718 2707 722
rect 2781 718 2785 722
rect 2865 718 2869 722
rect 2935 718 2939 722
rect 2436 706 2440 710
rect 2464 706 2468 710
rect 2796 708 2800 712
rect 2824 708 2828 712
rect 1616 663 1620 667
rect 1756 664 1760 668
rect 374 592 378 596
rect 467 592 471 596
rect 554 592 558 596
rect 1756 594 1760 598
rect 1616 585 1620 589
rect 1606 570 1610 574
rect 1766 553 1770 557
rect 1606 542 1610 546
rect 198 519 202 523
rect 285 519 289 523
rect 378 519 382 523
rect 590 521 594 525
rect 683 521 687 525
rect 770 521 774 525
rect 1766 525 1770 529
rect 1756 510 1760 514
rect 1616 501 1620 505
rect 92 380 96 384
rect 170 380 174 384
rect 254 380 258 384
rect 324 380 328 384
rect 421 382 425 386
rect 499 382 503 386
rect 583 382 587 386
rect 1616 431 1620 435
rect 2063 448 2067 452
rect 1756 432 1760 436
rect 2150 448 2154 452
rect 2243 448 2247 452
rect 2455 450 2459 454
rect 2548 450 2552 454
rect 2635 450 2639 454
rect 653 382 657 386
rect 748 385 752 389
rect 826 385 830 389
rect 910 385 914 389
rect 980 385 984 389
rect 185 370 189 374
rect 213 370 217 374
rect 514 372 518 376
rect 542 372 546 376
rect 841 375 845 379
rect 869 375 873 379
rect 1453 344 1457 348
rect 91 234 95 238
rect 169 234 173 238
rect 253 234 257 238
rect 323 234 327 238
rect 420 236 424 240
rect 498 236 502 240
rect 582 236 586 240
rect 1748 308 1752 312
rect 1957 309 1961 313
rect 2035 309 2039 313
rect 2119 309 2123 313
rect 2189 309 2193 313
rect 2286 311 2290 315
rect 2364 311 2368 315
rect 2448 311 2452 315
rect 2518 311 2522 315
rect 2613 314 2617 318
rect 2691 314 2695 318
rect 2775 314 2779 318
rect 2845 314 2849 318
rect 2050 299 2054 303
rect 2078 299 2082 303
rect 2379 301 2383 305
rect 2407 301 2411 305
rect 2706 304 2710 308
rect 2734 304 2738 308
rect 652 236 656 240
rect 747 239 751 243
rect 825 239 829 243
rect 909 239 913 243
rect 979 239 983 243
rect 184 224 188 228
rect 212 224 216 228
rect 513 226 517 230
rect 541 226 545 230
rect 840 229 844 233
rect 868 229 872 233
rect 1748 238 1752 242
rect 1455 191 1459 195
rect 1758 197 1762 201
rect 1457 165 1461 169
rect 1758 169 1762 173
rect 1956 163 1960 167
rect 2034 163 2038 167
rect 2118 163 2122 167
rect 2188 163 2192 167
rect 2285 165 2289 169
rect 2363 165 2367 169
rect 2447 165 2451 169
rect 2517 165 2521 169
rect 2612 168 2616 172
rect 2690 168 2694 172
rect 2774 168 2778 172
rect 2844 168 2848 172
rect 1748 154 1752 158
rect 2049 153 2053 157
rect 2077 153 2081 157
rect 2378 155 2382 159
rect 2406 155 2410 159
rect 2705 158 2709 162
rect 2733 158 2737 162
rect 385 86 389 90
rect 478 86 482 90
rect 565 86 569 90
rect 1748 76 1752 80
rect 2250 15 2254 19
rect 2343 15 2347 19
rect 2430 15 2434 19
<< nsubstratencontact >>
rect 1694 1052 1698 1056
rect 1694 1038 1698 1042
rect 1215 1027 1219 1031
rect 1269 1027 1273 1031
rect 1325 1027 1329 1031
rect 1379 1027 1383 1031
rect 1674 1023 1678 1027
rect 1694 1024 1698 1028
rect 1674 1009 1678 1013
rect 1674 995 1678 999
rect 1694 987 1698 991
rect 187 965 191 969
rect 274 965 278 969
rect 367 965 371 969
rect 579 967 583 971
rect 672 967 676 971
rect 759 967 763 971
rect 81 946 85 950
rect 95 946 99 950
rect 109 946 113 950
rect 192 946 196 950
rect 276 946 280 950
rect 313 946 317 950
rect 327 946 331 950
rect 341 946 345 950
rect 410 948 414 952
rect 424 948 428 952
rect 438 948 442 952
rect 521 948 525 952
rect 605 948 609 952
rect 642 948 646 952
rect 656 948 660 952
rect 670 948 674 952
rect 737 951 741 955
rect 751 951 755 955
rect 765 951 769 955
rect 848 951 852 955
rect 932 951 936 955
rect 969 951 973 955
rect 983 951 987 955
rect 997 951 1001 955
rect 1219 900 1223 904
rect 1273 900 1277 904
rect 1329 900 1333 904
rect 1383 900 1387 904
rect 1544 902 1548 906
rect 2453 926 2457 930
rect 1674 912 1678 916
rect 1694 903 1698 907
rect 1421 886 1425 890
rect 1215 882 1219 886
rect 1269 882 1273 886
rect 1325 882 1329 886
rect 1379 882 1383 886
rect 1824 913 1828 917
rect 2813 928 2817 932
rect 202 816 206 820
rect 531 818 535 822
rect 858 821 862 825
rect 1674 828 1678 832
rect 80 800 84 804
rect 94 800 98 804
rect 108 800 112 804
rect 191 800 195 804
rect 275 800 279 804
rect 312 800 316 804
rect 326 800 330 804
rect 340 800 344 804
rect 409 802 413 806
rect 423 802 427 806
rect 437 802 441 806
rect 520 802 524 806
rect 604 802 608 806
rect 641 802 645 806
rect 655 802 659 806
rect 669 802 673 806
rect 736 805 740 809
rect 750 805 754 809
rect 764 805 768 809
rect 847 805 851 809
rect 931 805 935 809
rect 968 805 972 809
rect 982 805 986 809
rect 996 805 1000 809
rect 1694 820 1698 824
rect 1694 806 1698 810
rect 1674 791 1678 795
rect 1694 792 1698 796
rect 1219 755 1223 759
rect 1273 755 1277 759
rect 1329 755 1333 759
rect 1383 755 1387 759
rect 1422 757 1426 761
rect 2314 796 2318 800
rect 2328 796 2332 800
rect 2342 796 2346 800
rect 2379 796 2383 800
rect 2463 796 2467 800
rect 2546 796 2550 800
rect 2560 796 2564 800
rect 2574 796 2578 800
rect 2674 798 2678 802
rect 2688 798 2692 802
rect 2702 798 2706 802
rect 2739 798 2743 802
rect 2823 798 2827 802
rect 2906 798 2910 802
rect 2920 798 2924 802
rect 2934 798 2938 802
rect 1987 784 1991 788
rect 2001 784 2005 788
rect 2015 784 2019 788
rect 1674 777 1678 781
rect 1674 763 1678 767
rect 1421 746 1425 750
rect 1214 740 1218 744
rect 1268 740 1272 744
rect 1324 740 1328 744
rect 1378 740 1382 744
rect 2098 784 2102 788
rect 2182 784 2186 788
rect 2219 784 2223 788
rect 2233 784 2237 788
rect 2247 784 2251 788
rect 2343 776 2347 780
rect 2357 776 2361 780
rect 2371 776 2375 780
rect 2454 776 2458 780
rect 2538 776 2542 780
rect 2575 776 2579 780
rect 2589 776 2593 780
rect 2603 776 2607 780
rect 2703 778 2707 782
rect 2717 778 2721 782
rect 2731 778 2735 782
rect 1696 692 1700 696
rect 2814 778 2818 782
rect 2898 778 2902 782
rect 2935 778 2939 782
rect 2949 778 2953 782
rect 2963 778 2967 782
rect 201 670 205 674
rect 530 672 534 676
rect 857 675 861 679
rect 1696 678 1700 682
rect 374 652 378 656
rect 467 652 471 656
rect 554 652 558 656
rect 1676 663 1680 667
rect 1696 664 1700 668
rect 1676 649 1680 653
rect 1676 635 1680 639
rect 2108 654 2112 658
rect 2464 646 2468 650
rect 2824 648 2828 652
rect 1696 627 1700 631
rect 1218 613 1222 617
rect 1272 613 1276 617
rect 1328 613 1332 617
rect 1382 613 1386 617
rect 1546 542 1550 546
rect 1676 552 1680 556
rect 1696 543 1700 547
rect 1236 516 1240 520
rect 1290 516 1294 520
rect 1346 516 1350 520
rect 1400 516 1404 520
rect 1826 553 1830 557
rect 198 459 202 463
rect 285 459 289 463
rect 378 459 382 463
rect 590 461 594 465
rect 683 461 687 465
rect 770 461 774 465
rect 1676 468 1680 472
rect 1696 460 1700 464
rect 92 440 96 444
rect 106 440 110 444
rect 120 440 124 444
rect 203 440 207 444
rect 287 440 291 444
rect 324 440 328 444
rect 338 440 342 444
rect 352 440 356 444
rect 421 442 425 446
rect 435 442 439 446
rect 449 442 453 446
rect 532 442 536 446
rect 616 442 620 446
rect 653 442 657 446
rect 667 442 671 446
rect 681 442 685 446
rect 748 445 752 449
rect 762 445 766 449
rect 776 445 780 449
rect 859 445 863 449
rect 943 445 947 449
rect 980 445 984 449
rect 994 445 998 449
rect 1008 445 1012 449
rect 1696 446 1700 450
rect 1676 431 1680 435
rect 1696 432 1700 436
rect 1676 417 1680 421
rect 1676 403 1680 407
rect 1240 389 1244 393
rect 1294 389 1298 393
rect 1350 389 1354 393
rect 1404 389 1408 393
rect 2063 388 2067 392
rect 2150 388 2154 392
rect 2243 388 2247 392
rect 2455 390 2459 394
rect 2548 390 2552 394
rect 2635 390 2639 394
rect 1234 371 1238 375
rect 1288 371 1292 375
rect 1344 371 1348 375
rect 1398 371 1402 375
rect 1957 369 1961 373
rect 1971 369 1975 373
rect 1985 369 1989 373
rect 213 310 217 314
rect 542 312 546 316
rect 869 315 873 319
rect 1688 336 1692 340
rect 1688 322 1692 326
rect 91 294 95 298
rect 105 294 109 298
rect 119 294 123 298
rect 202 294 206 298
rect 286 294 290 298
rect 323 294 327 298
rect 337 294 341 298
rect 351 294 355 298
rect 420 296 424 300
rect 434 296 438 300
rect 448 296 452 300
rect 531 296 535 300
rect 615 296 619 300
rect 652 296 656 300
rect 666 296 670 300
rect 680 296 684 300
rect 747 299 751 303
rect 761 299 765 303
rect 775 299 779 303
rect 858 299 862 303
rect 942 299 946 303
rect 979 299 983 303
rect 993 299 997 303
rect 1007 299 1011 303
rect 1453 284 1457 288
rect 2068 369 2072 373
rect 2152 369 2156 373
rect 2189 369 2193 373
rect 2203 369 2207 373
rect 2217 369 2221 373
rect 2286 371 2290 375
rect 2300 371 2304 375
rect 2314 371 2318 375
rect 1688 308 1692 312
rect 2397 371 2401 375
rect 2481 371 2485 375
rect 2518 371 2522 375
rect 2532 371 2536 375
rect 2546 371 2550 375
rect 2613 374 2617 378
rect 2627 374 2631 378
rect 2641 374 2645 378
rect 2724 374 2728 378
rect 2808 374 2812 378
rect 2845 374 2849 378
rect 2859 374 2863 378
rect 2873 374 2877 378
rect 1688 271 1692 275
rect 1455 251 1459 255
rect 1238 244 1242 248
rect 1292 244 1296 248
rect 1348 244 1352 248
rect 1402 244 1406 248
rect 1235 229 1239 233
rect 1289 229 1293 233
rect 1345 229 1349 233
rect 1399 229 1403 233
rect 2078 239 2082 243
rect 2407 241 2411 245
rect 2734 244 2738 248
rect 1956 223 1960 227
rect 1970 223 1974 227
rect 1984 223 1988 227
rect 1688 187 1692 191
rect 212 164 216 168
rect 541 166 545 170
rect 868 169 872 173
rect 385 146 389 150
rect 478 146 482 150
rect 565 146 569 150
rect 1818 197 1822 201
rect 2067 223 2071 227
rect 2151 223 2155 227
rect 2188 223 2192 227
rect 2202 223 2206 227
rect 2216 223 2220 227
rect 2285 225 2289 229
rect 2299 225 2303 229
rect 2313 225 2317 229
rect 2396 225 2400 229
rect 2480 225 2484 229
rect 2517 225 2521 229
rect 2531 225 2535 229
rect 2545 225 2549 229
rect 2612 228 2616 232
rect 2626 228 2630 232
rect 2640 228 2644 232
rect 2723 228 2727 232
rect 2807 228 2811 232
rect 2844 228 2848 232
rect 2858 228 2862 232
rect 2872 228 2876 232
rect 1239 102 1243 106
rect 1293 102 1297 106
rect 1349 102 1353 106
rect 1403 102 1407 106
rect 1457 105 1461 109
rect 1688 104 1692 108
rect 1688 90 1692 94
rect 2077 93 2081 97
rect 2406 95 2410 99
rect 2733 98 2737 102
rect 1688 76 1692 80
rect 2250 75 2254 79
rect 2343 75 2347 79
rect 2430 75 2434 79
<< psubstratepdiff >>
rect 578 1031 584 1032
rect 186 1029 192 1030
rect 186 1025 187 1029
rect 191 1025 192 1029
rect 186 1024 192 1025
rect 273 1029 279 1030
rect 273 1025 274 1029
rect 278 1025 279 1029
rect 273 1024 279 1025
rect 366 1029 372 1030
rect 366 1025 367 1029
rect 371 1025 372 1029
rect 578 1027 579 1031
rect 583 1027 584 1031
rect 578 1026 584 1027
rect 671 1031 677 1032
rect 671 1027 672 1031
rect 676 1027 677 1031
rect 366 1024 372 1025
rect 671 1026 677 1027
rect 758 1031 764 1032
rect 758 1027 759 1031
rect 763 1027 764 1031
rect 758 1026 764 1027
rect 1613 1027 1619 1028
rect 1613 1023 1614 1027
rect 1618 1023 1619 1027
rect 1613 1022 1619 1023
rect 1753 1028 1759 1029
rect 1753 1024 1754 1028
rect 1758 1024 1759 1028
rect 1753 1023 1759 1024
rect 80 890 86 891
rect 80 886 81 890
rect 85 886 86 890
rect 80 885 86 886
rect 158 890 164 891
rect 158 886 159 890
rect 163 886 164 890
rect 158 885 164 886
rect 242 890 248 891
rect 242 886 243 890
rect 247 886 248 890
rect 242 885 248 886
rect 409 892 415 893
rect 312 890 318 891
rect 312 886 313 890
rect 317 886 318 890
rect 312 885 318 886
rect 409 888 410 892
rect 414 888 415 892
rect 409 887 415 888
rect 487 892 493 893
rect 487 888 488 892
rect 492 888 493 892
rect 487 887 493 888
rect 571 892 577 893
rect 571 888 572 892
rect 576 888 577 892
rect 571 887 577 888
rect 1753 958 1759 959
rect 1753 954 1754 958
rect 1758 954 1759 958
rect 1753 953 1759 954
rect 1613 949 1619 950
rect 1613 945 1614 949
rect 1618 945 1619 949
rect 1613 944 1619 945
rect 736 895 742 896
rect 641 892 647 893
rect 641 888 642 892
rect 646 888 647 892
rect 641 887 647 888
rect 736 891 737 895
rect 741 891 742 895
rect 736 890 742 891
rect 814 895 820 896
rect 814 891 815 895
rect 819 891 820 895
rect 814 890 820 891
rect 898 895 904 896
rect 898 891 899 895
rect 903 891 904 895
rect 898 890 904 891
rect 1603 934 1609 935
rect 1603 930 1604 934
rect 1608 930 1609 934
rect 1603 906 1609 930
rect 1763 917 1769 918
rect 1763 913 1764 917
rect 1768 913 1769 917
rect 1603 902 1604 906
rect 1608 902 1609 906
rect 1603 901 1609 902
rect 968 895 974 896
rect 968 891 969 895
rect 973 891 974 895
rect 968 890 974 891
rect 829 885 863 886
rect 502 882 536 883
rect 173 880 207 881
rect 173 876 174 880
rect 178 876 202 880
rect 206 876 207 880
rect 502 878 503 882
rect 507 878 531 882
rect 535 878 536 882
rect 829 881 830 885
rect 834 881 858 885
rect 862 881 863 885
rect 829 880 863 881
rect 502 877 536 878
rect 173 875 207 876
rect 1763 889 1769 913
rect 1763 885 1764 889
rect 1768 885 1769 889
rect 1763 884 1769 885
rect 1753 874 1759 875
rect 1753 870 1754 874
rect 1758 870 1759 874
rect 1753 869 1759 870
rect 2452 870 2486 871
rect 1613 865 1619 866
rect 1613 861 1614 865
rect 1618 861 1619 865
rect 1613 860 1619 861
rect 2452 866 2453 870
rect 2457 866 2481 870
rect 2485 866 2486 870
rect 2812 872 2846 873
rect 2812 868 2813 872
rect 2817 868 2841 872
rect 2845 868 2846 872
rect 2812 867 2846 868
rect 2452 865 2486 866
rect 2341 860 2347 861
rect 2341 856 2342 860
rect 2346 856 2347 860
rect 2341 855 2347 856
rect 1420 830 1426 831
rect 1420 826 1421 830
rect 1425 826 1426 830
rect 1420 825 1426 826
rect 2411 860 2417 861
rect 2411 856 2412 860
rect 2416 856 2417 860
rect 2411 855 2417 856
rect 2495 860 2501 861
rect 2495 856 2496 860
rect 2500 856 2501 860
rect 2495 855 2501 856
rect 2573 860 2579 861
rect 2573 856 2574 860
rect 2578 856 2579 860
rect 2701 862 2707 863
rect 2701 858 2702 862
rect 2706 858 2707 862
rect 2701 857 2707 858
rect 2573 855 2579 856
rect 1421 821 1427 822
rect 1421 817 1422 821
rect 1426 817 1427 821
rect 1421 816 1427 817
rect 79 744 85 745
rect 79 740 80 744
rect 84 740 85 744
rect 79 739 85 740
rect 157 744 163 745
rect 157 740 158 744
rect 162 740 163 744
rect 157 739 163 740
rect 241 744 247 745
rect 241 740 242 744
rect 246 740 247 744
rect 241 739 247 740
rect 408 746 414 747
rect 311 744 317 745
rect 311 740 312 744
rect 316 740 317 744
rect 311 739 317 740
rect 408 742 409 746
rect 413 742 414 746
rect 408 741 414 742
rect 486 746 492 747
rect 486 742 487 746
rect 491 742 492 746
rect 486 741 492 742
rect 570 746 576 747
rect 570 742 571 746
rect 575 742 576 746
rect 570 741 576 742
rect 1613 795 1619 796
rect 1613 791 1614 795
rect 1618 791 1619 795
rect 1613 790 1619 791
rect 735 749 741 750
rect 640 746 646 747
rect 640 742 641 746
rect 645 742 646 746
rect 640 741 646 742
rect 735 745 736 749
rect 740 745 741 749
rect 735 744 741 745
rect 813 749 819 750
rect 813 745 814 749
rect 818 745 819 749
rect 813 744 819 745
rect 897 749 903 750
rect 897 745 898 749
rect 902 745 903 749
rect 897 744 903 745
rect 1753 796 1759 797
rect 1753 792 1754 796
rect 1758 792 1759 796
rect 2771 862 2777 863
rect 2771 858 2772 862
rect 2776 858 2777 862
rect 2771 857 2777 858
rect 2855 862 2861 863
rect 2855 858 2856 862
rect 2860 858 2861 862
rect 2855 857 2861 858
rect 2933 862 2939 863
rect 2933 858 2934 862
rect 2938 858 2939 862
rect 2933 857 2939 858
rect 1753 791 1759 792
rect 967 749 973 750
rect 967 745 968 749
rect 972 745 973 749
rect 967 744 973 745
rect 828 739 862 740
rect 501 736 535 737
rect 172 734 206 735
rect 172 730 173 734
rect 177 730 201 734
rect 205 730 206 734
rect 501 732 502 736
rect 506 732 530 736
rect 534 732 535 736
rect 828 735 829 739
rect 833 735 857 739
rect 861 735 862 739
rect 828 734 862 735
rect 501 731 535 732
rect 172 729 206 730
rect 1986 728 1992 729
rect 1986 724 1987 728
rect 1991 724 1992 728
rect 1986 723 1992 724
rect 2064 728 2070 729
rect 2064 724 2065 728
rect 2069 724 2070 728
rect 2064 723 2070 724
rect 2148 728 2154 729
rect 2148 724 2149 728
rect 2153 724 2154 728
rect 2148 723 2154 724
rect 2218 728 2224 729
rect 2218 724 2219 728
rect 2223 724 2224 728
rect 2218 723 2224 724
rect 1420 690 1426 691
rect 1420 686 1421 690
rect 1425 686 1426 690
rect 1420 685 1426 686
rect 2342 720 2348 721
rect 2079 718 2113 719
rect 2079 714 2080 718
rect 2084 714 2108 718
rect 2112 714 2113 718
rect 2342 716 2343 720
rect 2347 716 2348 720
rect 2342 715 2348 716
rect 2420 720 2426 721
rect 2420 716 2421 720
rect 2425 716 2426 720
rect 2420 715 2426 716
rect 2504 720 2510 721
rect 2504 716 2505 720
rect 2509 716 2510 720
rect 2504 715 2510 716
rect 2702 722 2708 723
rect 2574 720 2580 721
rect 2574 716 2575 720
rect 2579 716 2580 720
rect 2574 715 2580 716
rect 2702 718 2703 722
rect 2707 718 2708 722
rect 2702 717 2708 718
rect 2780 722 2786 723
rect 2780 718 2781 722
rect 2785 718 2786 722
rect 2780 717 2786 718
rect 2864 722 2870 723
rect 2864 718 2865 722
rect 2869 718 2870 722
rect 2864 717 2870 718
rect 2934 722 2940 723
rect 2934 718 2935 722
rect 2939 718 2940 722
rect 2934 717 2940 718
rect 2079 713 2113 714
rect 2795 712 2829 713
rect 2435 710 2469 711
rect 2435 706 2436 710
rect 2440 706 2464 710
rect 2468 706 2469 710
rect 2795 708 2796 712
rect 2800 708 2824 712
rect 2828 708 2829 712
rect 2795 707 2829 708
rect 2435 705 2469 706
rect 1615 667 1621 668
rect 1615 663 1616 667
rect 1620 663 1621 667
rect 1615 662 1621 663
rect 1755 668 1761 669
rect 1755 664 1756 668
rect 1760 664 1761 668
rect 1755 663 1761 664
rect 373 596 379 597
rect 373 592 374 596
rect 378 592 379 596
rect 373 591 379 592
rect 466 596 472 597
rect 466 592 467 596
rect 471 592 472 596
rect 466 591 472 592
rect 553 596 559 597
rect 553 592 554 596
rect 558 592 559 596
rect 553 591 559 592
rect 1755 598 1761 599
rect 1755 594 1756 598
rect 1760 594 1761 598
rect 1755 593 1761 594
rect 1615 589 1621 590
rect 1615 585 1616 589
rect 1620 585 1621 589
rect 1615 584 1621 585
rect 1605 574 1611 575
rect 1605 570 1606 574
rect 1610 570 1611 574
rect 1605 546 1611 570
rect 1765 557 1771 558
rect 1765 553 1766 557
rect 1770 553 1771 557
rect 1605 542 1606 546
rect 1610 542 1611 546
rect 1605 541 1611 542
rect 589 525 595 526
rect 197 523 203 524
rect 197 519 198 523
rect 202 519 203 523
rect 197 518 203 519
rect 284 523 290 524
rect 284 519 285 523
rect 289 519 290 523
rect 284 518 290 519
rect 377 523 383 524
rect 377 519 378 523
rect 382 519 383 523
rect 589 521 590 525
rect 594 521 595 525
rect 589 520 595 521
rect 682 525 688 526
rect 682 521 683 525
rect 687 521 688 525
rect 377 518 383 519
rect 682 520 688 521
rect 769 525 775 526
rect 769 521 770 525
rect 774 521 775 525
rect 769 520 775 521
rect 1765 529 1771 553
rect 1765 525 1766 529
rect 1770 525 1771 529
rect 1765 524 1771 525
rect 1755 514 1761 515
rect 1755 510 1756 514
rect 1760 510 1761 514
rect 1755 509 1761 510
rect 1615 505 1621 506
rect 1615 501 1616 505
rect 1620 501 1621 505
rect 1615 500 1621 501
rect 91 384 97 385
rect 91 380 92 384
rect 96 380 97 384
rect 91 379 97 380
rect 169 384 175 385
rect 169 380 170 384
rect 174 380 175 384
rect 169 379 175 380
rect 253 384 259 385
rect 253 380 254 384
rect 258 380 259 384
rect 253 379 259 380
rect 420 386 426 387
rect 323 384 329 385
rect 323 380 324 384
rect 328 380 329 384
rect 323 379 329 380
rect 420 382 421 386
rect 425 382 426 386
rect 420 381 426 382
rect 498 386 504 387
rect 498 382 499 386
rect 503 382 504 386
rect 498 381 504 382
rect 582 386 588 387
rect 582 382 583 386
rect 587 382 588 386
rect 582 381 588 382
rect 2454 454 2460 455
rect 1615 435 1621 436
rect 1615 431 1616 435
rect 1620 431 1621 435
rect 1615 430 1621 431
rect 2062 452 2068 453
rect 2062 448 2063 452
rect 2067 448 2068 452
rect 2062 447 2068 448
rect 1755 436 1761 437
rect 1755 432 1756 436
rect 1760 432 1761 436
rect 2149 452 2155 453
rect 2149 448 2150 452
rect 2154 448 2155 452
rect 2149 447 2155 448
rect 2242 452 2248 453
rect 2242 448 2243 452
rect 2247 448 2248 452
rect 2454 450 2455 454
rect 2459 450 2460 454
rect 2454 449 2460 450
rect 2547 454 2553 455
rect 2547 450 2548 454
rect 2552 450 2553 454
rect 2242 447 2248 448
rect 2547 449 2553 450
rect 2634 454 2640 455
rect 2634 450 2635 454
rect 2639 450 2640 454
rect 2634 449 2640 450
rect 1755 431 1761 432
rect 747 389 753 390
rect 652 386 658 387
rect 652 382 653 386
rect 657 382 658 386
rect 652 381 658 382
rect 747 385 748 389
rect 752 385 753 389
rect 747 384 753 385
rect 825 389 831 390
rect 825 385 826 389
rect 830 385 831 389
rect 825 384 831 385
rect 909 389 915 390
rect 909 385 910 389
rect 914 385 915 389
rect 909 384 915 385
rect 979 389 985 390
rect 979 385 980 389
rect 984 385 985 389
rect 979 384 985 385
rect 840 379 874 380
rect 513 376 547 377
rect 184 374 218 375
rect 184 370 185 374
rect 189 370 213 374
rect 217 370 218 374
rect 513 372 514 376
rect 518 372 542 376
rect 546 372 547 376
rect 840 375 841 379
rect 845 375 869 379
rect 873 375 874 379
rect 840 374 874 375
rect 513 371 547 372
rect 184 369 218 370
rect 1452 348 1458 349
rect 1452 344 1453 348
rect 1457 344 1458 348
rect 1452 343 1458 344
rect 90 238 96 239
rect 90 234 91 238
rect 95 234 96 238
rect 90 233 96 234
rect 168 238 174 239
rect 168 234 169 238
rect 173 234 174 238
rect 168 233 174 234
rect 252 238 258 239
rect 252 234 253 238
rect 257 234 258 238
rect 252 233 258 234
rect 419 240 425 241
rect 322 238 328 239
rect 322 234 323 238
rect 327 234 328 238
rect 322 233 328 234
rect 419 236 420 240
rect 424 236 425 240
rect 419 235 425 236
rect 497 240 503 241
rect 497 236 498 240
rect 502 236 503 240
rect 497 235 503 236
rect 581 240 587 241
rect 581 236 582 240
rect 586 236 587 240
rect 581 235 587 236
rect 1956 313 1962 314
rect 1747 312 1753 313
rect 1747 308 1748 312
rect 1752 308 1753 312
rect 1956 309 1957 313
rect 1961 309 1962 313
rect 1956 308 1962 309
rect 2034 313 2040 314
rect 2034 309 2035 313
rect 2039 309 2040 313
rect 2034 308 2040 309
rect 1747 307 1753 308
rect 2118 313 2124 314
rect 2118 309 2119 313
rect 2123 309 2124 313
rect 2118 308 2124 309
rect 2285 315 2291 316
rect 2188 313 2194 314
rect 2188 309 2189 313
rect 2193 309 2194 313
rect 2188 308 2194 309
rect 2285 311 2286 315
rect 2290 311 2291 315
rect 2285 310 2291 311
rect 2363 315 2369 316
rect 2363 311 2364 315
rect 2368 311 2369 315
rect 2363 310 2369 311
rect 2447 315 2453 316
rect 2447 311 2448 315
rect 2452 311 2453 315
rect 2447 310 2453 311
rect 2612 318 2618 319
rect 2517 315 2523 316
rect 2517 311 2518 315
rect 2522 311 2523 315
rect 2517 310 2523 311
rect 2612 314 2613 318
rect 2617 314 2618 318
rect 2612 313 2618 314
rect 2690 318 2696 319
rect 2690 314 2691 318
rect 2695 314 2696 318
rect 2690 313 2696 314
rect 2774 318 2780 319
rect 2774 314 2775 318
rect 2779 314 2780 318
rect 2774 313 2780 314
rect 2844 318 2850 319
rect 2844 314 2845 318
rect 2849 314 2850 318
rect 2844 313 2850 314
rect 2705 308 2739 309
rect 2378 305 2412 306
rect 2049 303 2083 304
rect 2049 299 2050 303
rect 2054 299 2078 303
rect 2082 299 2083 303
rect 2378 301 2379 305
rect 2383 301 2407 305
rect 2411 301 2412 305
rect 2705 304 2706 308
rect 2710 304 2734 308
rect 2738 304 2739 308
rect 2705 303 2739 304
rect 2378 300 2412 301
rect 2049 298 2083 299
rect 746 243 752 244
rect 651 240 657 241
rect 651 236 652 240
rect 656 236 657 240
rect 651 235 657 236
rect 746 239 747 243
rect 751 239 752 243
rect 746 238 752 239
rect 824 243 830 244
rect 824 239 825 243
rect 829 239 830 243
rect 824 238 830 239
rect 908 243 914 244
rect 908 239 909 243
rect 913 239 914 243
rect 908 238 914 239
rect 978 243 984 244
rect 978 239 979 243
rect 983 239 984 243
rect 978 238 984 239
rect 839 233 873 234
rect 512 230 546 231
rect 183 228 217 229
rect 183 224 184 228
rect 188 224 212 228
rect 216 224 217 228
rect 512 226 513 230
rect 517 226 541 230
rect 545 226 546 230
rect 839 229 840 233
rect 844 229 868 233
rect 872 229 873 233
rect 839 228 873 229
rect 512 225 546 226
rect 183 223 217 224
rect 1747 242 1753 243
rect 1747 238 1748 242
rect 1752 238 1753 242
rect 1747 237 1753 238
rect 1454 195 1460 196
rect 1454 191 1455 195
rect 1459 191 1460 195
rect 1757 201 1763 202
rect 1757 197 1758 201
rect 1762 197 1763 201
rect 1454 190 1460 191
rect 1456 169 1462 170
rect 1456 165 1457 169
rect 1461 165 1462 169
rect 1456 164 1462 165
rect 1757 173 1763 197
rect 1757 169 1758 173
rect 1762 169 1763 173
rect 1757 168 1763 169
rect 1955 167 1961 168
rect 1955 163 1956 167
rect 1960 163 1961 167
rect 1955 162 1961 163
rect 2033 167 2039 168
rect 2033 163 2034 167
rect 2038 163 2039 167
rect 2033 162 2039 163
rect 2117 167 2123 168
rect 2117 163 2118 167
rect 2122 163 2123 167
rect 2117 162 2123 163
rect 2284 169 2290 170
rect 2187 167 2193 168
rect 2187 163 2188 167
rect 2192 163 2193 167
rect 2187 162 2193 163
rect 2284 165 2285 169
rect 2289 165 2290 169
rect 2284 164 2290 165
rect 2362 169 2368 170
rect 2362 165 2363 169
rect 2367 165 2368 169
rect 2362 164 2368 165
rect 2446 169 2452 170
rect 2446 165 2447 169
rect 2451 165 2452 169
rect 2446 164 2452 165
rect 2611 172 2617 173
rect 2516 169 2522 170
rect 2516 165 2517 169
rect 2521 165 2522 169
rect 2516 164 2522 165
rect 2611 168 2612 172
rect 2616 168 2617 172
rect 2611 167 2617 168
rect 2689 172 2695 173
rect 2689 168 2690 172
rect 2694 168 2695 172
rect 2689 167 2695 168
rect 2773 172 2779 173
rect 2773 168 2774 172
rect 2778 168 2779 172
rect 2773 167 2779 168
rect 2843 172 2849 173
rect 2843 168 2844 172
rect 2848 168 2849 172
rect 2843 167 2849 168
rect 2704 162 2738 163
rect 2377 159 2411 160
rect 1747 158 1753 159
rect 1747 154 1748 158
rect 1752 154 1753 158
rect 2048 157 2082 158
rect 1747 153 1753 154
rect 2048 153 2049 157
rect 2053 153 2077 157
rect 2081 153 2082 157
rect 2377 155 2378 159
rect 2382 155 2406 159
rect 2410 155 2411 159
rect 2704 158 2705 162
rect 2709 158 2733 162
rect 2737 158 2738 162
rect 2704 157 2738 158
rect 2377 154 2411 155
rect 2048 152 2082 153
rect 384 90 390 91
rect 384 86 385 90
rect 389 86 390 90
rect 384 85 390 86
rect 477 90 483 91
rect 477 86 478 90
rect 482 86 483 90
rect 477 85 483 86
rect 564 90 570 91
rect 564 86 565 90
rect 569 86 570 90
rect 564 85 570 86
rect 1747 80 1753 81
rect 1747 76 1748 80
rect 1752 76 1753 80
rect 1747 75 1753 76
rect 2249 19 2255 20
rect 2249 15 2250 19
rect 2254 15 2255 19
rect 2249 14 2255 15
rect 2342 19 2348 20
rect 2342 15 2343 19
rect 2347 15 2348 19
rect 2342 14 2348 15
rect 2429 19 2435 20
rect 2429 15 2430 19
rect 2434 15 2435 19
rect 2429 14 2435 15
<< nsubstratendiff >>
rect 1693 1056 1699 1057
rect 1693 1052 1694 1056
rect 1698 1052 1699 1056
rect 1693 1042 1699 1052
rect 1693 1038 1694 1042
rect 1698 1038 1699 1042
rect 1693 1028 1699 1038
rect 1673 1027 1679 1028
rect 1673 1023 1674 1027
rect 1678 1023 1679 1027
rect 1693 1024 1694 1028
rect 1698 1024 1699 1028
rect 1693 1023 1699 1024
rect 1673 1013 1679 1023
rect 186 969 192 970
rect 273 969 279 970
rect 578 971 584 972
rect 1673 1009 1674 1013
rect 1678 1009 1679 1013
rect 671 971 677 972
rect 758 971 764 972
rect 1673 999 1679 1009
rect 1673 995 1674 999
rect 1678 995 1679 999
rect 1673 994 1679 995
rect 1693 991 1699 992
rect 1693 987 1694 991
rect 1698 987 1699 991
rect 1693 986 1699 987
rect 366 969 372 970
rect 186 965 187 969
rect 191 965 192 969
rect 186 964 192 965
rect 273 965 274 969
rect 278 965 279 969
rect 273 964 279 965
rect 366 965 367 969
rect 371 965 372 969
rect 578 967 579 971
rect 583 967 584 971
rect 578 966 584 967
rect 671 967 672 971
rect 676 967 677 971
rect 671 966 677 967
rect 758 967 759 971
rect 763 967 764 971
rect 758 966 764 967
rect 366 964 372 965
rect 409 952 443 953
rect 80 950 114 951
rect 80 946 81 950
rect 85 946 95 950
rect 99 946 109 950
rect 113 946 114 950
rect 191 950 197 951
rect 80 945 114 946
rect 191 946 192 950
rect 196 946 197 950
rect 275 950 281 951
rect 191 945 197 946
rect 275 946 276 950
rect 280 946 281 950
rect 312 950 346 951
rect 275 945 281 946
rect 312 946 313 950
rect 317 946 327 950
rect 331 946 341 950
rect 345 946 346 950
rect 409 948 410 952
rect 414 948 424 952
rect 428 948 438 952
rect 442 948 443 952
rect 520 952 526 953
rect 409 947 443 948
rect 312 945 346 946
rect 520 948 521 952
rect 525 948 526 952
rect 604 952 610 953
rect 520 947 526 948
rect 604 948 605 952
rect 609 948 610 952
rect 641 952 675 953
rect 604 947 610 948
rect 641 948 642 952
rect 646 948 656 952
rect 660 948 670 952
rect 674 948 675 952
rect 736 951 737 955
rect 741 951 751 955
rect 755 951 765 955
rect 769 951 770 955
rect 847 955 853 956
rect 736 950 770 951
rect 641 947 675 948
rect 847 951 848 955
rect 852 951 853 955
rect 931 955 937 956
rect 847 950 853 951
rect 931 951 932 955
rect 936 951 937 955
rect 968 955 1002 956
rect 931 950 937 951
rect 968 951 969 955
rect 973 951 983 955
rect 987 951 997 955
rect 1001 951 1002 955
rect 968 950 1002 951
rect 1543 906 1549 907
rect 1543 902 1544 906
rect 1548 902 1549 906
rect 1543 901 1549 902
rect 2452 930 2458 931
rect 2452 926 2453 930
rect 2457 926 2458 930
rect 2452 925 2458 926
rect 1673 916 1679 917
rect 1673 912 1674 916
rect 1678 912 1679 916
rect 1673 911 1679 912
rect 1693 907 1699 908
rect 1693 903 1694 907
rect 1698 903 1699 907
rect 1693 902 1699 903
rect 1420 890 1426 891
rect 1420 886 1421 890
rect 1425 886 1426 890
rect 1420 885 1426 886
rect 1823 917 1829 918
rect 1823 913 1824 917
rect 1828 913 1829 917
rect 1823 912 1829 913
rect 2812 932 2818 933
rect 2812 928 2813 932
rect 2817 928 2818 932
rect 2812 927 2818 928
rect 201 820 207 821
rect 857 825 863 826
rect 530 822 536 823
rect 201 816 202 820
rect 206 816 207 820
rect 530 818 531 822
rect 535 818 536 822
rect 857 821 858 825
rect 862 821 863 825
rect 1673 832 1679 833
rect 1673 828 1674 832
rect 1678 828 1679 832
rect 1673 827 1679 828
rect 1693 824 1699 825
rect 857 820 863 821
rect 530 817 536 818
rect 201 815 207 816
rect 735 809 769 810
rect 408 806 442 807
rect 79 804 113 805
rect 79 800 80 804
rect 84 800 94 804
rect 98 800 108 804
rect 112 800 113 804
rect 190 804 196 805
rect 79 799 113 800
rect 190 800 191 804
rect 195 800 196 804
rect 274 804 280 805
rect 190 799 196 800
rect 274 800 275 804
rect 279 800 280 804
rect 311 804 345 805
rect 274 799 280 800
rect 311 800 312 804
rect 316 800 326 804
rect 330 800 340 804
rect 344 800 345 804
rect 408 802 409 806
rect 413 802 423 806
rect 427 802 437 806
rect 441 802 442 806
rect 519 806 525 807
rect 408 801 442 802
rect 311 799 345 800
rect 519 802 520 806
rect 524 802 525 806
rect 603 806 609 807
rect 519 801 525 802
rect 603 802 604 806
rect 608 802 609 806
rect 640 806 674 807
rect 603 801 609 802
rect 640 802 641 806
rect 645 802 655 806
rect 659 802 669 806
rect 673 802 674 806
rect 735 805 736 809
rect 740 805 750 809
rect 754 805 764 809
rect 768 805 769 809
rect 846 809 852 810
rect 735 804 769 805
rect 640 801 674 802
rect 846 805 847 809
rect 851 805 852 809
rect 930 809 936 810
rect 846 804 852 805
rect 930 805 931 809
rect 935 805 936 809
rect 967 809 1001 810
rect 930 804 936 805
rect 967 805 968 809
rect 972 805 982 809
rect 986 805 996 809
rect 1000 805 1001 809
rect 967 804 1001 805
rect 1693 820 1694 824
rect 1698 820 1699 824
rect 1693 810 1699 820
rect 1693 806 1694 810
rect 1698 806 1699 810
rect 1693 796 1699 806
rect 2313 800 2347 801
rect 1673 795 1679 796
rect 1673 791 1674 795
rect 1678 791 1679 795
rect 1693 792 1694 796
rect 1698 792 1699 796
rect 1693 791 1699 792
rect 1421 761 1427 762
rect 1421 757 1422 761
rect 1426 757 1427 761
rect 1421 756 1427 757
rect 1673 781 1679 791
rect 2313 796 2314 800
rect 2318 796 2328 800
rect 2332 796 2342 800
rect 2346 796 2347 800
rect 2378 800 2384 801
rect 2313 795 2347 796
rect 2378 796 2379 800
rect 2383 796 2384 800
rect 2462 800 2468 801
rect 2378 795 2384 796
rect 2462 796 2463 800
rect 2467 796 2468 800
rect 2673 802 2707 803
rect 2545 800 2579 801
rect 2462 795 2468 796
rect 2545 796 2546 800
rect 2550 796 2560 800
rect 2564 796 2574 800
rect 2578 796 2579 800
rect 2673 798 2674 802
rect 2678 798 2688 802
rect 2692 798 2702 802
rect 2706 798 2707 802
rect 2738 802 2744 803
rect 2673 797 2707 798
rect 2738 798 2739 802
rect 2743 798 2744 802
rect 2822 802 2828 803
rect 2738 797 2744 798
rect 2822 798 2823 802
rect 2827 798 2828 802
rect 2905 802 2939 803
rect 2822 797 2828 798
rect 2905 798 2906 802
rect 2910 798 2920 802
rect 2924 798 2934 802
rect 2938 798 2939 802
rect 2905 797 2939 798
rect 2545 795 2579 796
rect 1986 788 2020 789
rect 1986 784 1987 788
rect 1991 784 2001 788
rect 2005 784 2015 788
rect 2019 784 2020 788
rect 2097 788 2103 789
rect 1986 783 2020 784
rect 1673 777 1674 781
rect 1678 777 1679 781
rect 1673 767 1679 777
rect 1673 763 1674 767
rect 1678 763 1679 767
rect 1673 762 1679 763
rect 1420 750 1426 751
rect 1420 746 1421 750
rect 1425 746 1426 750
rect 1420 745 1426 746
rect 2097 784 2098 788
rect 2102 784 2103 788
rect 2181 788 2187 789
rect 2097 783 2103 784
rect 2181 784 2182 788
rect 2186 784 2187 788
rect 2218 788 2252 789
rect 2181 783 2187 784
rect 2218 784 2219 788
rect 2223 784 2233 788
rect 2237 784 2247 788
rect 2251 784 2252 788
rect 2218 783 2252 784
rect 2702 782 2736 783
rect 2342 780 2376 781
rect 2342 776 2343 780
rect 2347 776 2357 780
rect 2361 776 2371 780
rect 2375 776 2376 780
rect 2453 780 2459 781
rect 2342 775 2376 776
rect 2453 776 2454 780
rect 2458 776 2459 780
rect 2537 780 2543 781
rect 2453 775 2459 776
rect 2537 776 2538 780
rect 2542 776 2543 780
rect 2574 780 2608 781
rect 2537 775 2543 776
rect 2574 776 2575 780
rect 2579 776 2589 780
rect 2593 776 2603 780
rect 2607 776 2608 780
rect 2702 778 2703 782
rect 2707 778 2717 782
rect 2721 778 2731 782
rect 2735 778 2736 782
rect 2813 782 2819 783
rect 2702 777 2736 778
rect 2574 775 2608 776
rect 200 674 206 675
rect 1695 696 1701 697
rect 1695 692 1696 696
rect 1700 692 1701 696
rect 1695 682 1701 692
rect 2813 778 2814 782
rect 2818 778 2819 782
rect 2897 782 2903 783
rect 2813 777 2819 778
rect 2897 778 2898 782
rect 2902 778 2903 782
rect 2934 782 2968 783
rect 2897 777 2903 778
rect 2934 778 2935 782
rect 2939 778 2949 782
rect 2953 778 2963 782
rect 2967 778 2968 782
rect 2934 777 2968 778
rect 856 679 862 680
rect 529 676 535 677
rect 200 670 201 674
rect 205 670 206 674
rect 529 672 530 676
rect 534 672 535 676
rect 856 675 857 679
rect 861 675 862 679
rect 856 674 862 675
rect 1695 678 1696 682
rect 1700 678 1701 682
rect 529 671 535 672
rect 200 669 206 670
rect 373 656 379 657
rect 373 652 374 656
rect 378 652 379 656
rect 466 656 472 657
rect 466 652 467 656
rect 471 652 472 656
rect 553 656 559 657
rect 553 652 554 656
rect 558 652 559 656
rect 373 651 379 652
rect 466 651 472 652
rect 553 651 559 652
rect 1695 668 1701 678
rect 1675 667 1681 668
rect 1675 663 1676 667
rect 1680 663 1681 667
rect 1695 664 1696 668
rect 1700 664 1701 668
rect 1695 663 1701 664
rect 1675 653 1681 663
rect 1675 649 1676 653
rect 1680 649 1681 653
rect 1675 639 1681 649
rect 1675 635 1676 639
rect 1680 635 1681 639
rect 2107 658 2113 659
rect 2107 654 2108 658
rect 2112 654 2113 658
rect 2107 653 2113 654
rect 2463 650 2469 651
rect 2823 652 2829 653
rect 2463 646 2464 650
rect 2468 646 2469 650
rect 2823 648 2824 652
rect 2828 648 2829 652
rect 2823 647 2829 648
rect 2463 645 2469 646
rect 1675 634 1681 635
rect 1695 631 1701 632
rect 1695 627 1696 631
rect 1700 627 1701 631
rect 1695 626 1701 627
rect 1545 546 1551 547
rect 1545 542 1546 546
rect 1550 542 1551 546
rect 1545 541 1551 542
rect 1675 556 1681 557
rect 1675 552 1676 556
rect 1680 552 1681 556
rect 1675 551 1681 552
rect 1695 547 1701 548
rect 1695 543 1696 547
rect 1700 543 1701 547
rect 1695 542 1701 543
rect 1825 557 1831 558
rect 1825 553 1826 557
rect 1830 553 1831 557
rect 1825 552 1831 553
rect 197 463 203 464
rect 284 463 290 464
rect 589 465 595 466
rect 682 465 688 466
rect 769 465 775 466
rect 377 463 383 464
rect 197 459 198 463
rect 202 459 203 463
rect 197 458 203 459
rect 284 459 285 463
rect 289 459 290 463
rect 284 458 290 459
rect 377 459 378 463
rect 382 459 383 463
rect 589 461 590 465
rect 594 461 595 465
rect 589 460 595 461
rect 682 461 683 465
rect 687 461 688 465
rect 682 460 688 461
rect 769 461 770 465
rect 774 461 775 465
rect 1675 472 1681 473
rect 1675 468 1676 472
rect 1680 468 1681 472
rect 1675 467 1681 468
rect 1695 464 1701 465
rect 769 460 775 461
rect 377 458 383 459
rect 1695 460 1696 464
rect 1700 460 1701 464
rect 420 446 454 447
rect 91 444 125 445
rect 91 440 92 444
rect 96 440 106 444
rect 110 440 120 444
rect 124 440 125 444
rect 202 444 208 445
rect 91 439 125 440
rect 202 440 203 444
rect 207 440 208 444
rect 286 444 292 445
rect 202 439 208 440
rect 286 440 287 444
rect 291 440 292 444
rect 323 444 357 445
rect 286 439 292 440
rect 323 440 324 444
rect 328 440 338 444
rect 342 440 352 444
rect 356 440 357 444
rect 420 442 421 446
rect 425 442 435 446
rect 439 442 449 446
rect 453 442 454 446
rect 531 446 537 447
rect 420 441 454 442
rect 323 439 357 440
rect 531 442 532 446
rect 536 442 537 446
rect 615 446 621 447
rect 531 441 537 442
rect 615 442 616 446
rect 620 442 621 446
rect 652 446 686 447
rect 615 441 621 442
rect 652 442 653 446
rect 657 442 667 446
rect 671 442 681 446
rect 685 442 686 446
rect 747 445 748 449
rect 752 445 762 449
rect 766 445 776 449
rect 780 445 781 449
rect 858 449 864 450
rect 747 444 781 445
rect 652 441 686 442
rect 858 445 859 449
rect 863 445 864 449
rect 942 449 948 450
rect 858 444 864 445
rect 942 445 943 449
rect 947 445 948 449
rect 979 449 1013 450
rect 942 444 948 445
rect 979 445 980 449
rect 984 445 994 449
rect 998 445 1008 449
rect 1012 445 1013 449
rect 1695 450 1701 460
rect 1695 446 1696 450
rect 1700 446 1701 450
rect 979 444 1013 445
rect 1695 436 1701 446
rect 1675 435 1681 436
rect 1675 431 1676 435
rect 1680 431 1681 435
rect 1695 432 1696 436
rect 1700 432 1701 436
rect 1695 431 1701 432
rect 1675 421 1681 431
rect 1675 417 1676 421
rect 1680 417 1681 421
rect 1675 407 1681 417
rect 1675 403 1676 407
rect 1680 403 1681 407
rect 1675 402 1681 403
rect 2062 392 2068 393
rect 2149 392 2155 393
rect 2454 394 2460 395
rect 2547 394 2553 395
rect 2634 394 2640 395
rect 2242 392 2248 393
rect 2062 388 2063 392
rect 2067 388 2068 392
rect 2062 387 2068 388
rect 2149 388 2150 392
rect 2154 388 2155 392
rect 2149 387 2155 388
rect 2242 388 2243 392
rect 2247 388 2248 392
rect 2454 390 2455 394
rect 2459 390 2460 394
rect 2454 389 2460 390
rect 2547 390 2548 394
rect 2552 390 2553 394
rect 2547 389 2553 390
rect 2634 390 2635 394
rect 2639 390 2640 394
rect 2634 389 2640 390
rect 2242 387 2248 388
rect 2285 375 2319 376
rect 1956 373 1990 374
rect 1956 369 1957 373
rect 1961 369 1971 373
rect 1975 369 1985 373
rect 1989 369 1990 373
rect 2067 373 2073 374
rect 1956 368 1990 369
rect 212 314 218 315
rect 868 319 874 320
rect 541 316 547 317
rect 212 310 213 314
rect 217 310 218 314
rect 541 312 542 316
rect 546 312 547 316
rect 868 315 869 319
rect 873 315 874 319
rect 1687 340 1693 341
rect 1687 336 1688 340
rect 1692 336 1693 340
rect 1687 326 1693 336
rect 868 314 874 315
rect 1687 322 1688 326
rect 1692 322 1693 326
rect 541 311 547 312
rect 212 309 218 310
rect 746 303 780 304
rect 419 300 453 301
rect 90 298 124 299
rect 90 294 91 298
rect 95 294 105 298
rect 109 294 119 298
rect 123 294 124 298
rect 201 298 207 299
rect 90 293 124 294
rect 201 294 202 298
rect 206 294 207 298
rect 285 298 291 299
rect 201 293 207 294
rect 285 294 286 298
rect 290 294 291 298
rect 322 298 356 299
rect 285 293 291 294
rect 322 294 323 298
rect 327 294 337 298
rect 341 294 351 298
rect 355 294 356 298
rect 419 296 420 300
rect 424 296 434 300
rect 438 296 448 300
rect 452 296 453 300
rect 530 300 536 301
rect 419 295 453 296
rect 322 293 356 294
rect 530 296 531 300
rect 535 296 536 300
rect 614 300 620 301
rect 530 295 536 296
rect 614 296 615 300
rect 619 296 620 300
rect 651 300 685 301
rect 614 295 620 296
rect 651 296 652 300
rect 656 296 666 300
rect 670 296 680 300
rect 684 296 685 300
rect 746 299 747 303
rect 751 299 761 303
rect 765 299 775 303
rect 779 299 780 303
rect 857 303 863 304
rect 746 298 780 299
rect 651 295 685 296
rect 857 299 858 303
rect 862 299 863 303
rect 941 303 947 304
rect 857 298 863 299
rect 941 299 942 303
rect 946 299 947 303
rect 978 303 1012 304
rect 941 298 947 299
rect 978 299 979 303
rect 983 299 993 303
rect 997 299 1007 303
rect 1011 299 1012 303
rect 978 298 1012 299
rect 1452 288 1458 289
rect 1452 284 1453 288
rect 1457 284 1458 288
rect 1452 283 1458 284
rect 1687 312 1693 322
rect 2067 369 2068 373
rect 2072 369 2073 373
rect 2151 373 2157 374
rect 2067 368 2073 369
rect 2151 369 2152 373
rect 2156 369 2157 373
rect 2188 373 2222 374
rect 2151 368 2157 369
rect 2188 369 2189 373
rect 2193 369 2203 373
rect 2207 369 2217 373
rect 2221 369 2222 373
rect 2285 371 2286 375
rect 2290 371 2300 375
rect 2304 371 2314 375
rect 2318 371 2319 375
rect 2396 375 2402 376
rect 2285 370 2319 371
rect 2188 368 2222 369
rect 1687 308 1688 312
rect 1692 308 1693 312
rect 1687 307 1693 308
rect 2396 371 2397 375
rect 2401 371 2402 375
rect 2480 375 2486 376
rect 2396 370 2402 371
rect 2480 371 2481 375
rect 2485 371 2486 375
rect 2517 375 2551 376
rect 2480 370 2486 371
rect 2517 371 2518 375
rect 2522 371 2532 375
rect 2536 371 2546 375
rect 2550 371 2551 375
rect 2612 374 2613 378
rect 2617 374 2627 378
rect 2631 374 2641 378
rect 2645 374 2646 378
rect 2723 378 2729 379
rect 2612 373 2646 374
rect 2517 370 2551 371
rect 2723 374 2724 378
rect 2728 374 2729 378
rect 2807 378 2813 379
rect 2723 373 2729 374
rect 2807 374 2808 378
rect 2812 374 2813 378
rect 2844 378 2878 379
rect 2807 373 2813 374
rect 2844 374 2845 378
rect 2849 374 2859 378
rect 2863 374 2873 378
rect 2877 374 2878 378
rect 2844 373 2878 374
rect 1687 275 1693 276
rect 1687 271 1688 275
rect 1692 271 1693 275
rect 1687 270 1693 271
rect 1454 255 1460 256
rect 1454 251 1455 255
rect 1459 251 1460 255
rect 1454 250 1460 251
rect 2077 243 2083 244
rect 2733 248 2739 249
rect 2406 245 2412 246
rect 2077 239 2078 243
rect 2082 239 2083 243
rect 2406 241 2407 245
rect 2411 241 2412 245
rect 2733 244 2734 248
rect 2738 244 2739 248
rect 2733 243 2739 244
rect 2406 240 2412 241
rect 2077 238 2083 239
rect 2611 232 2645 233
rect 2284 229 2318 230
rect 1955 227 1989 228
rect 1955 223 1956 227
rect 1960 223 1970 227
rect 1974 223 1984 227
rect 1988 223 1989 227
rect 2066 227 2072 228
rect 1955 222 1989 223
rect 211 168 217 169
rect 1687 191 1693 192
rect 1687 187 1688 191
rect 1692 187 1693 191
rect 1687 186 1693 187
rect 867 173 873 174
rect 540 170 546 171
rect 211 164 212 168
rect 216 164 217 168
rect 540 166 541 170
rect 545 166 546 170
rect 867 169 868 173
rect 872 169 873 173
rect 867 168 873 169
rect 540 165 546 166
rect 211 163 217 164
rect 384 150 390 151
rect 384 146 385 150
rect 389 146 390 150
rect 477 150 483 151
rect 477 146 478 150
rect 482 146 483 150
rect 564 150 570 151
rect 564 146 565 150
rect 569 146 570 150
rect 384 145 390 146
rect 477 145 483 146
rect 564 145 570 146
rect 1817 201 1823 202
rect 1817 197 1818 201
rect 1822 197 1823 201
rect 1817 196 1823 197
rect 2066 223 2067 227
rect 2071 223 2072 227
rect 2150 227 2156 228
rect 2066 222 2072 223
rect 2150 223 2151 227
rect 2155 223 2156 227
rect 2187 227 2221 228
rect 2150 222 2156 223
rect 2187 223 2188 227
rect 2192 223 2202 227
rect 2206 223 2216 227
rect 2220 223 2221 227
rect 2284 225 2285 229
rect 2289 225 2299 229
rect 2303 225 2313 229
rect 2317 225 2318 229
rect 2395 229 2401 230
rect 2284 224 2318 225
rect 2187 222 2221 223
rect 2395 225 2396 229
rect 2400 225 2401 229
rect 2479 229 2485 230
rect 2395 224 2401 225
rect 2479 225 2480 229
rect 2484 225 2485 229
rect 2516 229 2550 230
rect 2479 224 2485 225
rect 2516 225 2517 229
rect 2521 225 2531 229
rect 2535 225 2545 229
rect 2549 225 2550 229
rect 2611 228 2612 232
rect 2616 228 2626 232
rect 2630 228 2640 232
rect 2644 228 2645 232
rect 2722 232 2728 233
rect 2611 227 2645 228
rect 2516 224 2550 225
rect 2722 228 2723 232
rect 2727 228 2728 232
rect 2806 232 2812 233
rect 2722 227 2728 228
rect 2806 228 2807 232
rect 2811 228 2812 232
rect 2843 232 2877 233
rect 2806 227 2812 228
rect 2843 228 2844 232
rect 2848 228 2858 232
rect 2862 228 2872 232
rect 2876 228 2877 232
rect 2843 227 2877 228
rect 1456 109 1462 110
rect 1456 105 1457 109
rect 1461 105 1462 109
rect 1456 104 1462 105
rect 1687 108 1693 109
rect 1687 104 1688 108
rect 1692 104 1693 108
rect 1687 94 1693 104
rect 1687 90 1688 94
rect 1692 90 1693 94
rect 2076 97 2082 98
rect 2732 102 2738 103
rect 2405 99 2411 100
rect 1687 80 1693 90
rect 2076 93 2077 97
rect 2081 93 2082 97
rect 2405 95 2406 99
rect 2410 95 2411 99
rect 2732 98 2733 102
rect 2737 98 2738 102
rect 2732 97 2738 98
rect 2405 94 2411 95
rect 2076 92 2082 93
rect 1687 76 1688 80
rect 1692 76 1693 80
rect 1687 75 1693 76
rect 2249 79 2255 80
rect 2249 75 2250 79
rect 2254 75 2255 79
rect 2342 79 2348 80
rect 2342 75 2343 79
rect 2347 75 2348 79
rect 2429 79 2435 80
rect 2429 75 2430 79
rect 2434 75 2435 79
rect 2249 74 2255 75
rect 2342 74 2348 75
rect 2429 74 2435 75
<< pad >>
rect 214 959 218 963
rect 225 453 229 457
rect 2090 382 2094 386
<< labels >>
rlabel metal1 845 675 845 675 2 vdd
rlabel m2contact 155 1009 155 1009 1 q0_M1
rlabel metal1 191 1001 191 1001 1 q0b2_M1
rlabel metal1 363 1008 363 1008 1 q0b0_n_M1
rlabel metal1 483 1014 483 1014 1 b2_M1
rlabel metal1 484 993 484 993 1 b1_M1
rlabel metal1 484 974 484 974 1 b0_M1
rlabel metal1 578 1012 578 1012 1 q1b0_M1
rlabel metal1 680 1019 680 1019 1 q1b1_M1
rlabel metal1 680 997 680 997 1 q1b1_n_M1
rlabel metal1 758 1008 758 1008 1 q1b2_M1
rlabel metal1 767 1008 767 1008 1 q1b2_n_M1
rlabel m2contact 794 1011 794 1011 1 q1_M1
rlabel metal1 983 919 983 919 1 zc1_n_3_M1
rlabel metal1 969 919 969 919 1 c1_3_M1
rlabel metal1 955 923 955 923 1 s_fa3_M1
rlabel metal1 932 941 932 941 1 cn_3_M1
rlabel metal1 871 923 871 923 1 so_3_M1
rlabel metal1 859 944 859 944 1 bn3_M1
rlabel ptransistor 855 928 855 928 1 an3_M1
rlabel metal1 758 923 758 923 1 co_n3_M1
rlabel metal1 745 903 745 903 1 co_3_M1
rlabel metal1 642 916 642 916 1 c1_2_M1
rlabel metal1 656 916 656 916 1 zc1_2_n_M1
rlabel ntransistor 621 903 621 903 1 son_2_M1
rlabel pdcontact 618 933 618 933 1 s_fa2_M1
rlabel metal1 606 916 606 916 1 cn2_M1
rlabel metal1 544 920 544 920 1 so_2_M1
rlabel polycontact 534 916 534 916 1 an_2_M1
rlabel polycontact 528 917 528 917 1 bn_2_M1
rlabel metal1 431 919 431 919 1 co_n2_M1
rlabel metal1 418 900 418 900 1 co_2_M1
rlabel metal1 327 914 327 914 1 zc1_n1_M1
rlabel metal1 313 914 313 914 1 c1_1_M1
rlabel ntransistor 292 901 292 901 1 a1_n_M1
rlabel ntransistor 208 902 208 902 1 an_1_M1
rlabel metal1 215 918 215 918 1 so_1_M1
rlabel metal1 102 918 102 918 1 co_n1_M1
rlabel metal1 89 898 89 898 1 co_1_M1
rlabel metal1 198 846 198 846 1 c_fa1_n_M1
rlabel metal1 206 846 206 846 1 c_fa1_M1
rlabel metal1 527 850 527 850 1 c_fa_n_M1
rlabel metal1 535 854 535 854 1 c_fa2_M1
rlabel metal1 854 853 854 853 1 c_fa3_n_M1
rlabel metal1 862 857 862 857 1 c_fa3_M1
rlabel metal1 982 773 982 773 1 zc1_6_n_M1
rlabel metal1 968 773 968 773 1 c1_6_M1
rlabel ntransistor 947 760 947 760 1 s_fa_6_n_M1
rlabel metal1 930 794 930 794 1 cn_6_M1
rlabel metal1 870 777 870 777 1 so_6_M1
rlabel ptransistor 854 782 854 782 1 an_6_M1
rlabel metal1 815 771 815 771 1 bn_6_M1
rlabel metal1 757 777 757 777 1 co_n_6_M1
rlabel metal1 744 757 744 757 1 co_6_M1
rlabel metal1 655 770 655 770 1 zc1_n_5_M1
rlabel metal1 641 770 641 770 1 c1_5_M1
rlabel metal1 603 790 603 790 1 cn_5_M1
rlabel ntransistor 620 757 620 757 1 s_fa5_n_M1
rlabel metal1 531 795 531 795 1 bn_5_M1
rlabel ptransistor 527 779 527 779 1 an_5_M1
rlabel metal1 543 774 543 774 1 so_5_M1
rlabel metal1 430 774 430 774 1 co_5__M1
rlabel metal1 326 768 326 768 1 zc1_4_M1
rlabel metal1 312 768 312 768 1 c1_4_M1
rlabel ntransistor 291 755 291 755 1 s_fa4_n_M1
rlabel metal1 274 788 274 788 1 cn_1_M1
rlabel metal1 191 787 191 787 1 bn4_M1
rlabel ptransistor 198 777 198 777 1 an4_M1
rlabel metal1 214 772 214 772 1 so_4_M1
rlabel metal1 101 772 101 772 1 co_n4_M1
rlabel metal1 88 752 88 752 1 co_4_M1
rlabel metal1 197 702 197 702 1 a5_n_M1
rlabel metal1 534 708 534 708 1 c_fa5_M1
rlabel metal1 526 704 526 704 1 c_fa5_n_M1
rlabel metal1 853 707 853 707 1 c_fa6_n_M1
rlabel metal1 861 711 861 711 1 c_fa6_M1
rlabel metal1 554 614 554 614 1 q2b0_M1
rlabel metal1 563 613 563 613 1 q2b0_n_M1
rlabel m2contact 591 612 591 612 1 q2_M1
rlabel metal1 466 614 466 614 1 q2b1_M1
rlabel metal1 475 614 475 614 1 q2b1_n_M1
rlabel metal1 396 603 396 603 1 q2b2_n_M1
rlabel metal1 374 602 374 602 1 q2b2_M1
rlabel metal1 183 1005 183 1005 1 q0b2_n_M1
rlabel metal1 278 1005 278 1005 1 q0b1_M1
rlabel metal1 587 998 587 998 1 q1b0_n_M1
rlabel metal1 270 1006 270 1006 1 q0b1_n_M1
rlabel metal1 370 1007 370 1007 1 a0_M1
rlabel m2contact 1106 990 1106 990 1 en_bar_D1
rlabel metal1 1177 997 1177 997 1 D_bar_D1
rlabel metal1 1224 995 1224 995 1 out_n1_D1
rlabel ndiffusion 1205 978 1205 978 1 n1_D1
rlabel ndiffusion 1261 978 1261 978 1 n2_D1
rlabel metal1 1279 991 1279 991 1 out_n2_D1
rlabel ndiffusion 1317 978 1317 978 1 n3_D1
rlabel ndiffusion 1371 978 1371 978 1 n4_D1
rlabel m2contact 1388 994 1388 994 1 q_l1_bar_D1
rlabel m2contact 1392 937 1392 937 1 q_bar_D1
rlabel ndiffusion 1375 953 1375 953 1 n10_D1
rlabel metal1 1283 940 1283 940 1 out_n8_D1
rlabel ndiffusion 1265 953 1265 953 1 n8_D1
rlabel metal1 1228 936 1228 936 1 out_n7_D1
rlabel ndiffusion 1209 953 1209 953 1 n7_D1
rlabel polycontact 1199 933 1199 933 1 q_l1_D1
rlabel metal1 1181 937 1181 937 1 n6_D1
rlabel ndiffusion 1321 953 1321 953 1 n9_D1
rlabel m2contact 1338 929 1338 929 1 q_D1
rlabel m2contact 1388 849 1388 849 1 q_l1_bar_D2
rlabel metal1 1181 792 1181 792 1 n6_D2
rlabel polycontact 1199 788 1199 788 1 q_l1_D2
rlabel ndiffusion 1209 808 1209 808 1 n7_D2
rlabel metal1 1228 791 1228 791 1 out_n7__D2
rlabel ndiffusion 1265 808 1265 808 1 n8_D2
rlabel metal1 1283 795 1283 795 1 out_n8_D2
rlabel ndiffusion 1321 808 1321 808 1 n9_D2
rlabel m2contact 1338 784 1338 784 1 q_D2
rlabel ndiffusion 1375 808 1375 808 1 n10_D2
rlabel m2contact 1392 792 1392 792 1 q_bar_D2
rlabel ndiffusion 1371 833 1371 833 1 n4_D2
rlabel ndiffusion 1317 833 1317 833 1 n3_D2
rlabel metal1 1279 846 1279 846 1 out_n2_D2
rlabel ndiffusion 1261 833 1261 833 1 n2_D2
rlabel metal1 1224 850 1224 850 1 out_n1_D2
rlabel ndiffusion 1205 833 1205 833 1 n1_D2
rlabel metal1 1177 852 1177 852 1 D_bar_D2
rlabel m2contact 1106 845 1106 845 1 en_bar_D2
rlabel metal1 1180 650 1180 650 1 n6_D3
rlabel polycontact 1198 646 1198 646 1 q_l1_D3
rlabel metal1 1227 649 1227 649 1 out_n7_D3
rlabel ndiffusion 1264 666 1264 666 1 n8_D3
rlabel m2contact 1337 642 1337 642 1 q_D3
rlabel metal1 1282 653 1282 653 1 out_n8_D3
rlabel ndiffusion 1320 666 1320 666 1 n9_D3
rlabel m2contact 1391 650 1391 650 1 q_bar_D3
rlabel m2contact 1387 707 1387 707 1 q_l1_bar_D3
rlabel ndiffusion 1370 691 1370 691 1 n4_D3
rlabel ndiffusion 1316 691 1316 691 1 n3_D3
rlabel metal1 1278 704 1278 704 1 out_n2_D3
rlabel ndiffusion 1260 691 1260 691 1 n2_D3
rlabel metal1 1223 708 1223 708 1 out_n1_D3
rlabel ndiffusion 1204 691 1204 691 1 n1_D3
rlabel metal1 1176 710 1176 710 1 D_bar_D3
rlabel m2contact 1105 703 1105 703 1 en_bar_D3
rlabel ndiffusion 1374 666 1374 666 1 n10
rlabel polycontact 1216 998 1216 998 1 en
rlabel polycontact 1424 853 1424 853 1 q_D1
rlabel polycontact 1437 854 1437 854 1 q_D1_n
rlabel polycontact 1425 793 1425 793 1 q_D2
rlabel polycontact 1438 793 1438 793 1 q_n_D2
rlabel polycontact 1425 714 1425 714 1 q_D3
rlabel polycontact 1437 714 1437 714 1 q_D3_n
rlabel metal2 1433 125 1433 125 7 q_D6
rlabel metal1 1203 139 1203 139 1 n6_D6
rlabel polycontact 1219 135 1219 135 1 q_l1_D6
rlabel metal1 1248 138 1248 138 1 out_n7_D6
rlabel ndiffusion 1229 155 1229 155 1 n7_D6
rlabel metal1 1303 142 1303 142 1 out_n8_D6
rlabel ndiffusion 1285 155 1285 155 1 n8_D6
rlabel m2contact 1358 131 1358 131 1 q_D6
rlabel ndiffusion 1341 155 1341 155 1 n9_D6
rlabel m2contact 1412 139 1412 139 1 q_bar_D6
rlabel ndiffusion 1395 155 1395 155 1 n10_D6
rlabel m2contact 1408 196 1408 196 1 q_l1_bar_D6
rlabel ndiffusion 1391 180 1391 180 1 n4_D6
rlabel ndiffusion 1337 180 1337 180 1 n3_D6
rlabel metal1 1299 193 1299 193 1 out_n2_D6
rlabel ndiffusion 1281 180 1281 180 1 n2_D6
rlabel ndiffusion 1225 180 1225 180 1 n1_D6
rlabel metal1 1244 197 1244 197 1 out_n1_D6
rlabel metal1 1197 199 1197 199 1 D_Bar_D6
rlabel m2contact 1126 192 1126 192 1 en_bar_D6
rlabel metal2 1431 274 1431 274 7 q_D5
rlabel metal1 1201 281 1201 281 1 n6_D5
rlabel polycontact 1218 277 1218 277 1 q_l1_D5
rlabel metal1 1247 280 1247 280 1 out_n7_D5
rlabel ndiffusion 1284 297 1284 297 1 n8_D5
rlabel metal1 1302 284 1302 284 1 out_n8_D5
rlabel m2contact 1357 273 1357 273 1 q_D5
rlabel ndiffusion 1340 297 1340 297 1 n9_D5
rlabel metal1 1411 289 1411 289 1 q_bar_D5
rlabel ndiffusion 1394 297 1394 297 1 n10_D5
rlabel metal1 1407 343 1407 343 1 q_l1_bar_D5
rlabel ndiffusion 1390 322 1390 322 1 n4_D5
rlabel ndiffusion 1336 322 1336 322 1 n3_D5
rlabel metal1 1298 335 1298 335 1 out_n2_D5
rlabel ndiffusion 1280 322 1280 322 1 n2_D5
rlabel metal1 1243 339 1243 339 1 out_n1_D5
rlabel metal1 1196 341 1196 341 1 D_bar_D5
rlabel m2contact 1125 334 1125 334 1 en_bar_D5
rlabel metal1 1245 484 1245 484 1 out_n1_D4
rlabel metal1 1202 426 1202 426 1 n6_D4
rlabel polycontact 1220 422 1220 422 1 q_l1_D4
rlabel metal1 1249 425 1249 425 1 out_n7_D4
rlabel metal1 1304 429 1304 429 1 out_n8_D4
rlabel ndiffusion 1286 442 1286 442 1 n8_D4
rlabel ndiffusion 1342 442 1342 442 1 n9_D4
rlabel m2contact 1359 418 1359 418 1 q_D4
rlabel m2contact 1413 426 1413 426 1 q_bar_D4
rlabel ndiffusion 1396 442 1396 442 1 n10_D4
rlabel m2contact 1407 482 1407 482 1 q_l1_bar_D4
rlabel ndiffusion 1392 467 1392 467 1 n4_D4
rlabel ndiffusion 1338 467 1338 467 1 n3_D4
rlabel metal1 1300 480 1300 480 1 out_n2_D4
rlabel ndiffusion 1282 467 1282 467 1 n2_D4
rlabel metal1 1198 486 1198 486 1 D_bar_D4
rlabel m2contact 1127 479 1127 479 1 en_bar_D4
rlabel m2contact 166 503 166 503 1 q0_M2
rlabel metal1 194 499 194 499 1 q0b2_n_M2
rlabel metal1 202 495 202 495 1 q0b2_M2
rlabel metal1 281 500 281 500 1 q0b1_n_M2
rlabel metal1 289 499 289 499 1 q0b1_M2
rlabel metal1 374 502 374 502 1 q0b0_n_M2
rlabel metal1 494 508 494 508 1 b2_M2
rlabel metal1 495 468 495 468 1 b0_M2
rlabel metal1 495 487 495 487 1 b1_M2
rlabel metal1 691 513 691 513 1 q1b1_M2
rlabel metal1 769 502 769 502 1 q1b2_M2
rlabel metal1 778 502 778 502 1 q1b2_n_M2
rlabel m2contact 805 505 805 505 1 q1_M2
rlabel metal1 994 413 994 413 1 zc1_n_3_M2
rlabel metal1 980 413 980 413 1 c1_3_M2
rlabel metal1 966 417 966 417 1 s_fa3_M2
rlabel ntransistor 959 400 959 400 1 s_fa3_n_M2
rlabel metal1 882 417 882 417 1 so_3_M2
rlabel metal1 769 417 769 417 1 co_n3_M2
rlabel metal1 756 397 756 397 1 co_3_M2
rlabel metal1 667 410 667 410 1 zc1_2_n_M2
rlabel metal1 653 410 653 410 1 c1_2_M2
rlabel pdcontact 629 427 629 427 1 s_fa2_M2
rlabel metal1 617 410 617 410 1 cn2_M2
rlabel ntransistor 632 397 632 397 1 son_2_M2
rlabel metal1 555 414 555 414 1 so_2_M2
rlabel polycontact 538 411 538 411 1 bn_2_M2
rlabel polycontact 547 411 547 411 1 an_2_M2
rlabel metal1 442 413 442 413 1 co_n2_M2
rlabel metal1 429 394 429 394 1 co_2_M2
rlabel metal1 338 408 338 408 1 zc1_n1_M2
rlabel metal1 324 408 324 408 1 c1_1_M2
rlabel ntransistor 303 395 303 395 1 a1_1_M2
rlabel metal1 226 412 226 412 1 so_1_M2
rlabel ntransistor 219 396 219 396 1 an_1_M2
rlabel metal1 214 433 214 433 1 bn_1_M1
rlabel metal1 100 392 100 392 1 co_1_M2
rlabel metal1 113 412 113 412 1 co_n1_M2
rlabel metal1 209 340 209 340 1 c_fa1_n_M2
rlabel metal1 217 340 217 340 1 c_fa1_M2
rlabel metal1 538 344 538 344 1 c_fa2_n_M2
rlabel metal1 546 348 546 348 1 c_fa2_M2
rlabel metal1 865 347 865 347 1 c_fa3_n_M2
rlabel metal1 873 351 873 351 1 c_fa3_M2
rlabel metal1 993 267 993 267 1 zc1_6_n_M2
rlabel metal1 979 267 979 267 1 c1_6_M2
rlabel ntransistor 958 254 958 254 1 s_fa_6_n_M2
rlabel metal1 941 288 941 288 1 cn_6_M2
rlabel metal1 881 271 881 271 1 so_6_M2
rlabel ptransistor 865 276 865 276 1 an_6_M2
rlabel metal1 826 265 826 265 1 bn_6_M2
rlabel metal1 768 271 768 271 1 co_n_6_M2
rlabel metal1 755 251 755 251 1 co_6_M2
rlabel ntransistor 631 251 631 251 1 s_fa_5_n_M2
rlabel metal1 542 289 542 289 1 bn_5_M2
rlabel ptransistor 538 273 538 273 1 an_5_M2
rlabel metal1 554 268 554 268 1 so_5_M2
rlabel metal1 337 262 337 262 1 zc1_4_M2
rlabel metal1 323 262 323 262 1 c1_4_M2
rlabel ntransistor 302 249 302 249 1 s_fa4_n_M2
rlabel metal1 285 282 285 282 1 cn_1_M2
rlabel metal1 202 281 202 281 1 bn4_M2
rlabel ptransistor 209 271 209 271 1 an4_M2
rlabel metal1 225 266 225 266 1 so_4_M2
rlabel metal1 112 266 112 266 1 co_n4_M2
rlabel metal1 99 246 99 246 1 co_4_M2
rlabel polycontact 208 199 208 199 1 a5_n_M2
rlabel metal1 537 198 537 198 1 c_fa5_n_M2
rlabel metal1 545 202 545 202 1 c_fa5_M2
rlabel metal1 864 201 864 201 1 c_fa6_n_M2
rlabel metal1 872 205 872 205 1 c_fa6_M2
rlabel metal1 407 97 407 97 1 q2b2_n_M2
rlabel metal1 385 96 385 96 1 q2b2_M2
rlabel metal1 477 108 477 108 1 q2b1_M2
rlabel metal1 486 108 486 108 1 q2b1_n_M2
rlabel m2contact 602 106 602 106 1 q2_M2
rlabel metal1 574 107 574 107 1 q2b0_n_M2
rlabel metal1 565 108 565 108 1 q2b0_M2
rlabel metal1 589 506 589 506 1 q1b0_M2
rlabel metal1 598 492 598 492 1 q1b0_n_M2
rlabel metal1 943 435 943 435 1 cn_3_M2
rlabel ptransistor 866 422 866 422 1 an3_M2
rlabel metal1 870 438 870 438 1 bn3_M2
rlabel metal1 441 268 441 268 1 co_5_M2
rlabel metal1 691 491 691 491 1 q1b1_n_M2
rlabel metal1 66 498 66 498 1 q0_M2
rlabel metal2 64 546 64 546 5 q1_M2
rlabel metal1 345 106 346 106 1 q2_M2
rlabel metal2 1431 419 1431 419 1 q_D4
rlabel polycontact 1469 320 1469 320 1 q_D4_n
rlabel polycontact 1471 219 1472 219 1 q_D5_n
rlabel polycontact 1473 141 1473 141 1 q_D6_n
rlabel metal1 1720 97 1720 97 7 n1_A1
rlabel metal1 1740 84 1740 84 7 n5_A1
rlabel metal1 1704 154 1704 154 7 b1_A1
rlabel metal1 1699 198 1699 198 7 bn_A1
rlabel metal1 1726 155 1726 155 7 b1n_A1
rlabel polycontact 1728 170 1728 170 7 a1_A1
rlabel metal1 1720 210 1720 210 7 xor1_A1
rlabel ndcontact 1736 181 1736 181 7 a1n_A1
rlabel metal1 1705 270 1705 270 7 n3_A1
rlabel metal1 1720 294 1720 294 7 s1_A1
rlabel metal1 1724 308 1724 308 7 c1_A1
rlabel metal1 1724 322 1724 322 7 zc1_n_A1
rlabel metal1 1728 453 1728 453 7 n9_n_A1
rlabel metal1 1748 440 1748 440 7 n9_A1
rlabel metal1 1711 510 1711 510 7 b2_A1
rlabel metal1 1734 511 1734 511 7 b2n_A1
rlabel metal1 1740 518 1740 518 7 a2_A1
rlabel ptransistor 1723 550 1723 550 7 a2n_A1
rlabel metal1 1728 566 1728 566 7 xor_2_A1
rlabel metal2 1708 586 1708 586 7 s2_A1
rlabel metal1 1711 627 1711 627 7 n6_A1
rlabel metal1 1728 650 1728 650 7 s3_A1
rlabel ntransistor 1745 643 1745 643 7 n7_A1
rlabel metal1 1732 664 1732 664 7 n8_A1
rlabel metal1 1732 678 1732 678 7 zc2_n_A1
rlabel metal1 1628 659 1628 659 7 n10_A1
rlabel metal1 1648 646 1648 646 7 n10_nA1
rlabel m2contact 1713 391 1713 391 7 s2_A1
rlabel ntransistor 1632 540 1632 540 7 a3n_A1
rlabel polycontact 1640 573 1640 573 7 a3_A1
rlabel metal1 1648 533 1648 533 7 xor_3_A1
rlabel polycontact 1645 542 1645 542 7 a3n_A1
rlabel metal1 1645 557 1645 557 7 b3n_A1
rlabel metal1 1664 589 1664 589 7 b3_A1
rlabel m2contact 1582 542 1582 542 7 c3_A1
rlabel metal1 1578 550 1578 550 7 cout3_n_A1
rlabel metal1 1798 549 1798 549 7 cout2_n_A1
rlabel metal1 1795 557 1795 557 7 c2_A1
rlabel ntransistor 1631 456 1631 456 7 n11_A1
rlabel metal1 1648 449 1648 449 7 s4_a1
rlabel metal1 1664 477 1664 477 7 n12_A1
rlabel metal2 1668 497 1668 497 7 c2_A1
rlabel metal1 1644 435 1644 435 7 n13_A1
rlabel metal1 1644 421 1644 421 7 zc3_n_A1
rlabel metal1 1790 193 1790 193 7 cout_n_A1
rlabel metal1 1786 201 1786 201 7 s2_A1
rlabel metal1 1769 81 1769 81 7 co_A1
rlabel metal1 1772 112 1772 112 7 n2_A1
rlabel polycontact 1778 145 1778 145 7 son_A1
rlabel polycontact 1788 139 1788 139 7 con_A1
rlabel metal1 1785 153 1785 153 7 so_A1
rlabel metal1 1789 121 1789 121 7 b_A1
rlabel polycontact 1785 97 1785 97 7 a_A1
rlabel metal1 1642 781 1642 781 7 zc5_n_A1
rlabel metal1 1642 795 1642 795 7 n21_A1
rlabel ntransistor 1629 816 1629 816 7 n19_A1
rlabel metal1 1646 809 1646 809 7 s6_A1
rlabel metal1 1662 837 1662 837 7 n20_A1
rlabel metal2 1666 857 1666 857 7 c4_A1
rlabel ntransistor 1630 900 1630 900 7 a5n_A1
rlabel polycontact 1638 933 1638 933 7 a5_A1
rlabel metal1 1646 893 1646 893 7 xor_5_A1
rlabel metal1 1643 917 1643 917 7 b5n_A1
rlabel metal1 1662 949 1662 949 7 b5_A1
rlabel metal1 1626 1019 1626 1019 7 n18_A1
rlabel metal2 1711 751 1711 751 7 c3_A1
rlabel metal1 1726 813 1726 813 7 n17n_A1
rlabel metal1 1746 800 1746 800 7 n17_A1
rlabel metal1 1709 870 1709 870 7 b4_A1
rlabel metal1 1732 871 1732 871 7 b4n_A1
rlabel metal1 1738 878 1738 878 7 a4_A1
rlabel ptransistor 1721 910 1721 910 7 a4n_A1
rlabel metal1 1726 926 1726 926 7 xor_4_A1
rlabel metal2 1706 946 1706 946 7 c3_A1
rlabel metal1 1709 987 1709 987 7 n14_A1
rlabel metal1 1726 1010 1726 1010 7 s5_A1
rlabel ntransistor 1743 1003 1743 1003 7 n15_A1
rlabel metal1 1730 1024 1730 1024 7 n16_A1
rlabel metal1 1730 1038 1730 1038 7 zc4_n_A1
rlabel metal1 1792 917 1792 917 7 c4_A1
rlabel metal1 1796 909 1796 909 7 cout4n_A1
rlabel metal1 1576 910 1576 910 7 cout5_n_A1
rlabel metal1 1646 1006 1646 1006 7 n18_nA1
rlabel metal2 1720 27 1720 27 7 a1_A1
rlabel metal2 1842 23 1842 23 7 b2_A1
rlabel metal1 1591 332 1591 332 7 a3_A1
rlabel metal1 1601 331 1601 331 7 b3_A1
rlabel metal2 1853 24 1853 24 7 a4_A1
rlabel metal2 1868 21 1868 21 7 b4_A1
rlabel metal2 1551 440 1551 440 7 b5_A1
rlabel metal2 1534 435 1534 435 3 a5_A1
rlabel polycontact 1723 286 1723 286 7 n4_A1
rlabel metal2 1534 1066 1534 1066 4 s1_A1
rlabel metal1 1875 1075 1875 1075 7 so_A1
rlabel metal2 1840 1082 1840 1082 5 s3_A1
rlabel metal1 1860 1081 1860 1081 7 s1_A1
rlabel metal2 1826 1084 1826 1084 5 s5_A1
rlabel metal2 1816 1084 1816 1084 5 s6_A1
rlabel m2contact 1603 1076 1603 1076 7 s4_A1
rlabel metal2 1810 24 1810 24 1 a_A1
rlabel polysilicon 1815 23 1815 23 1 b_A1
rlabel metal2 1829 25 1829 25 1 a2_A1
rlabel polycontact 947 920 947 920 1 s_fa3_n_M1
rlabel polycontact 197 915 197 915 1 bn_n_M1
rlabel metal1 614 284 614 284 1 cn_5_M2
rlabel metal1 652 264 652 264 1 c1_5_M2
rlabel metal1 666 264 666 264 1 zc1_n_5_M2
rlabel metal1 249 1030 249 1030 1 vss
rlabel metal1 183 952 183 952 1 vdd
rlabel metal2 1707 26 1707 26 1 b1_A1
rlabel metal1 2395 305 2395 305 2 vss
rlabel m2contact 2031 432 2031 432 1 q0_M3
rlabel metal1 2059 428 2059 428 1 q0b2_n_M3
rlabel metal1 2067 424 2067 424 1 q0b2_M3
rlabel metal1 2146 429 2146 429 1 q0b1_n_M3
rlabel metal1 2154 428 2154 428 1 q0b1_M3
rlabel metal1 2239 431 2239 431 1 q0b0_n_M3
rlabel metal1 2359 437 2359 437 1 b2_M3
rlabel metal1 2360 416 2360 416 1 b1_M3
rlabel metal1 2360 397 2360 397 1 b0_M3
rlabel metal1 2454 435 2454 435 1 q1b0_M3
rlabel metal1 2463 421 2463 421 1 q1b0_n_M3
rlabel metal1 2556 442 2556 442 1 q1b1_M3
rlabel metal1 2556 420 2556 420 1 q1b1_n_M3
rlabel metal1 2643 431 2643 431 1 q1b2_n_M3
rlabel metal1 2845 342 2845 342 1 c1_3_M3
rlabel metal1 2859 342 2859 342 1 zc1_n_3_M3
rlabel metal1 2831 346 2831 346 1 s_fa3_M3
rlabel polycontact 2823 343 2823 343 1 s_fa3_n_M3
rlabel metal1 2808 364 2808 364 1 cn_3_M3
rlabel metal1 2747 346 2747 346 1 so_3_M3
rlabel ptransistor 2731 351 2731 351 1 an3_M3
rlabel metal1 2735 367 2735 367 1 bn3_M3
rlabel metal1 2634 346 2634 346 1 co_n3_M3
rlabel metal1 2621 326 2621 326 1 co_3_M3
rlabel metal1 2532 339 2532 339 1 zc1_n2_M3
rlabel metal1 2518 339 2518 339 1 c1_2_M3
rlabel ntransistor 2497 326 2497 326 1 son_2_M3
rlabel pdcontact 2494 356 2494 356 1 s_fa2_M3
rlabel metal1 2482 339 2482 339 1 cn_2_M3
rlabel metal1 2420 343 2420 343 1 so_2_M3
rlabel polycontact 2412 340 2412 340 1 an_2_M3
rlabel metal1 2307 343 2307 343 1 co_n2_M3
rlabel metal1 2294 323 2294 323 1 co_2_M3
rlabel metal1 2203 337 2203 337 1 zc1_n1_M3
rlabel metal1 2189 337 2189 337 1 c1_1_M3
rlabel metal1 2175 341 2175 341 1 a1_M3
rlabel metal1 2091 341 2091 341 1 so_1_M3
rlabel ntransistor 2084 325 2084 325 1 an_1_M3
rlabel metal1 2079 362 2079 362 1 bn_1_M3
rlabel metal1 1978 341 1978 341 1 co_n1_M3
rlabel metal1 1965 321 1965 321 1 co_1_M3
rlabel metal1 2082 269 2082 269 1 c_fa1_M3
rlabel metal1 2403 273 2403 273 1 c_fa2_n_M3
rlabel metal1 2738 280 2738 280 1 c_fa3_M3
rlabel metal1 2844 196 2844 196 1 c1_6_M3
rlabel metal1 2858 196 2858 196 1 zc1_n_6_M3
rlabel metal1 2830 200 2830 200 1 a2_M3
rlabel ntransistor 2823 183 2823 183 1 s_fa6_n_M3
rlabel metal1 2806 217 2806 217 1 cn_6_M3
rlabel ptransistor 2730 205 2730 205 1 an_6_M3
rlabel metal1 1964 175 1964 175 1 co_4_M3
rlabel metal1 1977 195 1977 195 1 co_n4_M3
rlabel metal1 2067 210 2067 210 1 bn4_M3
rlabel ptransistor 2074 200 2074 200 1 an4_M3
rlabel metal1 2090 195 2090 195 1 so_4_M3
rlabel metal1 2150 211 2150 211 1 cn_4_M3
rlabel metal1 2174 195 2174 195 1 a4_M3
rlabel metal1 2188 191 2188 191 1 c1_4_M3
rlabel metal1 2202 191 2202 191 1 zc1_4_M3
rlabel metal1 2306 197 2306 197 1 co_5_n_M3
rlabel metal1 2293 177 2293 177 1 co_5_M3
rlabel metal1 2407 218 2407 218 1 bn_5_M3
rlabel ptransistor 2403 202 2403 202 1 an_5_M3
rlabel metal1 2419 197 2419 197 1 so_5_M3
rlabel metal1 2479 213 2479 213 1 cn_5_M3
rlabel metal1 2503 197 2503 197 1 a3_M3
rlabel metal1 2517 193 2517 193 1 c1_5_M3
rlabel metal1 2531 193 2531 193 1 zc1_n_5_M3
rlabel metal1 2633 200 2633 200 1 co_n_6_M3
rlabel metal1 2620 180 2620 180 1 co_6_M3
rlabel metal1 2691 194 2691 194 1 bn_6_M3
rlabel metal1 2737 134 2737 134 1 c_fa6_M3
rlabel metal1 2729 130 2729 130 1 c_fa6_n_M3
rlabel metal1 2410 131 2410 131 1 c_fa5_M3
rlabel metal1 2402 127 2402 127 1 c_fa5_n_M3
rlabel metal1 2081 129 2081 129 1 a5_M3
rlabel metal1 2250 25 2250 25 1 q2b2_M3
rlabel metal1 2272 26 2272 26 1 q2b2_n_M3
rlabel metal1 2342 37 2342 37 1 q2b1_M3
rlabel metal1 2351 37 2351 37 1 q2b1_n_M3
rlabel metal1 2430 37 2430 37 1 q2b0_M3
rlabel metal1 2439 36 2439 36 1 q2b0_n_M3
rlabel m2contact 2467 35 2467 35 1 q2_M3
rlabel metal1 2634 431 2634 431 1 q1b2_M3
rlabel polycontact 2402 340 2402 340 1 bn_2_M3
rlabel metal1 2074 269 2074 269 1 c_fa1_n_M3
rlabel polycontact 2730 280 2730 280 1 c_fa3_n_M3
rlabel metal1 2746 200 2746 200 1 so_6_M3
rlabel m2contact 2489 435 2489 435 1 q1_M3
rlabel metal1 2246 430 2246 430 1 a0_M3
rlabel polycontact 2167 337 2167 337 1 a1_n_M3
rlabel polycontact 2166 192 2166 192 1 a4_n_M3
rlabel polycontact 2495 194 2495 194 1 a3_n_M3
rlabel polycontact 2073 128 2073 128 1 a5_n_M3
rlabel metal1 2461 898 2461 898 1 cout3_n_A2
rlabel m2contact 2453 894 2453 894 1 c3_A2
rlabel metal1 2813 896 2813 896 1 c5_A2
rlabel metal1 2821 900 2821 900 1 cout5_n_A2
rlabel metal1 2930 850 2930 850 1 n18_A2
rlabel metal1 2917 830 2917 830 1 n18_n_A2
rlabel polycontact 2844 838 2844 838 1 a5_A2
rlabel metal1 2828 833 2828 833 1 b5_n_A2
rlabel polycontact 2813 833 2813 833 1 a5_n_A2
rlabel metal1 2804 830 2804 830 1 xor_5_A2
rlabel m2contact 2770 810 2770 810 1 c4_A2
rlabel metal1 2748 814 2748 814 1 n20_A2
rlabel metal1 2720 830 2720 830 1 s6_A2
rlabel polycontact 2728 832 2728 832 1 n19_A2
rlabel metal1 2706 834 2706 834 1 n21_A2
rlabel metal1 2692 834 2692 834 1 zc5_n_A2
rlabel metal1 2570 848 2570 848 1 n10_A2
rlabel metal1 2557 828 2557 828 1 n1_n_A2
rlabel metal1 2468 831 2468 831 1 b3n_A2
rlabel polycontact 2453 831 2453 831 1 a3n_A2
rlabel metal1 2444 828 2444 828 1 xor_3_A2
rlabel metal2 2408 808 2408 808 1 c2_A2
rlabel metal1 2388 812 2388 812 1 n12_A2
rlabel metal1 2360 828 2360 828 1 s4_A2
rlabel ntransistor 2367 845 2367 845 1 n11_A2
rlabel metal1 2346 832 2346 832 1 n13_A2
rlabel metal1 2332 832 2332 832 1 zc3_n_A2
rlabel metal1 2949 746 2949 746 1 zc4_n_A2
rlabel metal1 2935 746 2935 746 1 n16_A2
rlabel metal1 2921 750 2921 750 1 s5_A2
rlabel metal1 2898 767 2898 767 1 n14_A2
rlabel metal2 2857 770 2857 770 1 c3_A2
rlabel metal1 2837 750 2837 750 1 xor_4_A2
rlabel ptransistor 2821 755 2821 755 1 a4n_A2
rlabel metal1 2782 744 2782 744 1 b4n_A2
rlabel metal1 2724 750 2724 750 1 n17_n_A2
rlabel metal1 2711 730 2711 730 1 n17_A2
rlabel metal2 2662 765 2662 765 1 c3_A2
rlabel metal1 2589 744 2589 744 1 zc2_n_A2
rlabel metal1 2575 744 2575 744 1 n8_A2
rlabel metal1 2561 748 2561 748 1 s3_A2
rlabel metal1 2538 765 2538 765 1 n6_A2
rlabel metal2 2497 768 2497 768 1 s2_A2
rlabel metal1 2477 748 2477 748 1 xor_2_A2
rlabel ptransistor 2461 753 2461 753 1 a2n_A2
rlabel metal1 2422 742 2422 742 1 b2n_A2
rlabel metal1 2351 728 2351 728 1 n9_A2
rlabel m2contact 2299 764 2299 764 1 s2_A2
rlabel metal1 2233 752 2233 752 1 zc1_n_A2
rlabel metal1 2219 752 2219 752 1 c1_A2
rlabel metal1 2205 756 2205 756 1 s1_A2
rlabel metal1 2181 771 2181 771 1 n3_A2
rlabel metal1 2121 756 2121 756 1 xor1_A2
rlabel metal1 2109 777 2109 777 1 bn_A2
rlabel ndcontact 2091 738 2091 738 1 a1n_A2
rlabel metal1 2066 750 2066 750 1 b1n_A2
rlabel metal1 1995 736 1995 736 1 n5_A2
rlabel ndcontact 1984 707 1984 707 1 co_A2
rlabel polycontact 1990 691 1990 691 1 con_A2
rlabel metal1 2023 704 2023 704 1 n2_A2
rlabel ntransistor 2038 700 2038 700 1 son_A2
rlabel polycontact 2050 688 2050 688 1 con_A2
rlabel metal1 2064 691 2064 691 1 so_A2
rlabel metal1 2112 690 2112 690 1 s2_A2
rlabel metal1 2468 682 2468 682 1 c2_A2
rlabel metal1 2460 678 2460 678 1 cout2_n_A2
rlabel metal1 2820 680 2820 680 1 cout4_n_A2
rlabel metal1 2828 684 2828 684 1 c4_A2
rlabel metal1 2104 686 2104 686 1 cout_n_A2
rlabel polycontact 2913 747 2913 747 1 n15_A2
rlabel polycontact 2553 745 2553 745 1 n7_A2
rlabel polycontact 2197 753 2197 753 1 n4_A2
rlabel metal1 2760 891 2760 891 1 s8_A2
rlabel metal1 2721 883 2721 883 1 n2_7_A2
rlabel polycontact 2688 889 2688 889 1 s7_n_A2
rlabel metal1 2680 896 2680 896 1 s7_A2
rlabel metal1 2008 754 2008 754 1 n1_A2
rlabel metal1 2364 745 2364 745 1 n9_n_A2
rlabel metal2 2982 889 2982 889 7 s8_A2
rlabel metal1 3004 984 3004 984 5 s7_A2
rlabel metal1 3006 1000 3006 1000 6 s4_A2
rlabel metal1 3001 1017 3001 1017 5 s1_A2
rlabel metal1 2955 626 2955 626 1 s3_A2
rlabel metal2 2983 753 2983 753 1 s5_A2
rlabel metal1 2957 589 2957 589 1 so_A2
rlabel metal2 2982 880 2982 880 1 s6_A2
rlabel metal2 1954 977 1954 977 1 c5_A2
rlabel metal1 2411 272 2411 272 1 c_fa2_M3
rlabel metal2 1939 964 1939 964 1 c5_A1
rlabel polycontact 1237 487 1237 487 1 en
rlabel ndiffusion 1235 297 1235 297 1 n7_D5
rlabel ndiffusion 1234 322 1234 322 1 n1_D5
rlabel ndiffusion 1235 441 1235 441 1 n7_D4
rlabel ndiffusion 1234 467 1234 467 1 n1_D4
rlabel ndiffusion 1217 666 1217 666 1 n7_D3
rlabel metal1 2729 912 2729 912 1 s8_n_A2
<< end >>
