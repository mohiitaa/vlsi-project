magic
tech scmos
timestamp 1521650470
<< pwell >>
rect -71 9 72 45
rect 84 9 202 45
rect 15 -17 63 9
<< nwell >>
rect -71 45 72 89
rect 84 45 202 89
rect 15 -24 63 -17
rect 11 -37 63 -24
rect 15 -61 63 -37
<< polysilicon >>
rect 21 79 23 83
rect -55 71 -49 72
rect -65 63 -63 68
rect -55 67 -54 71
rect -50 67 -49 71
rect -55 66 -49 67
rect -55 61 -53 66
rect -45 61 -43 66
rect 6 63 12 64
rect 6 59 7 63
rect 11 59 12 63
rect 6 58 12 59
rect -65 48 -63 51
rect -55 48 -53 51
rect -65 47 -59 48
rect -65 43 -64 47
rect -60 43 -59 47
rect -55 45 -51 48
rect -65 42 -59 43
rect -65 34 -63 42
rect -53 31 -51 45
rect -45 40 -43 51
rect 10 49 12 58
rect 57 79 59 83
rect 105 79 107 83
rect 37 70 39 74
rect 47 70 49 74
rect 90 63 96 64
rect 90 59 91 63
rect 95 59 96 63
rect 90 58 96 59
rect 21 49 23 52
rect 37 49 39 52
rect 47 49 49 52
rect 57 49 59 52
rect 10 47 23 49
rect 29 47 39 49
rect 43 48 49 49
rect -46 39 -40 40
rect 13 39 15 47
rect 29 43 31 47
rect 43 44 44 48
rect 48 44 49 48
rect 43 43 49 44
rect 53 48 59 49
rect 53 44 54 48
rect 58 44 59 48
rect 94 49 96 58
rect 141 79 143 83
rect 121 70 123 74
rect 131 70 133 74
rect 177 71 183 72
rect 167 63 169 68
rect 177 67 178 71
rect 182 67 183 71
rect 177 66 183 67
rect 105 49 107 52
rect 121 49 123 52
rect 131 49 133 52
rect 141 49 143 52
rect 177 61 179 66
rect 187 61 189 66
rect 94 47 107 49
rect 113 47 123 49
rect 127 48 133 49
rect 53 43 59 44
rect 22 42 31 43
rect -46 35 -45 39
rect -41 35 -40 39
rect -46 34 -40 35
rect -46 31 -44 34
rect -65 24 -63 28
rect 22 38 23 42
rect 27 38 31 42
rect 47 39 49 43
rect 22 37 31 38
rect 29 34 31 37
rect 39 34 41 39
rect 47 37 51 39
rect 49 34 51 37
rect 56 34 58 43
rect 97 39 99 47
rect 113 43 115 47
rect 127 44 128 48
rect 132 44 133 48
rect 127 43 133 44
rect 137 48 143 49
rect 137 44 138 48
rect 142 44 143 48
rect 137 43 143 44
rect 167 48 169 51
rect 177 48 179 51
rect 167 47 173 48
rect 167 43 168 47
rect 172 43 173 47
rect 177 45 181 48
rect 106 42 115 43
rect 13 27 15 30
rect 13 25 18 27
rect -53 17 -51 22
rect -46 17 -44 22
rect 16 17 18 25
rect 29 21 31 25
rect 39 17 41 25
rect 106 38 107 42
rect 111 38 115 42
rect 131 39 133 43
rect 106 37 115 38
rect 113 34 115 37
rect 123 34 125 39
rect 131 37 135 39
rect 133 34 135 37
rect 140 34 142 43
rect 167 42 173 43
rect 167 34 169 42
rect 97 27 99 30
rect 97 25 102 27
rect 49 17 51 22
rect 56 17 58 22
rect 16 15 41 17
rect 100 17 102 25
rect 113 21 115 25
rect 123 17 125 25
rect 179 31 181 45
rect 187 40 189 51
rect 186 39 192 40
rect 186 35 187 39
rect 191 35 192 39
rect 186 34 192 35
rect 186 31 188 34
rect 167 24 169 28
rect 133 17 135 22
rect 140 17 142 22
rect 100 15 125 17
rect 179 17 181 22
rect 186 17 188 22
rect 28 0 30 4
rect 38 0 40 4
rect 48 0 50 4
rect 28 -14 30 -6
rect 24 -15 30 -14
rect 38 -15 40 -6
rect 48 -15 50 -6
rect 24 -19 25 -15
rect 29 -19 30 -15
rect 44 -16 50 -15
rect 24 -20 30 -19
rect 28 -33 30 -20
rect 38 -22 40 -19
rect 44 -20 45 -16
rect 49 -20 50 -16
rect 44 -21 50 -20
rect 34 -23 40 -22
rect 34 -27 35 -23
rect 39 -27 40 -23
rect 34 -28 40 -27
rect 35 -33 37 -28
rect 48 -30 50 -21
rect 48 -46 50 -42
rect 28 -55 30 -51
rect 35 -55 37 -51
<< ndiffusion >>
rect -72 33 -65 34
rect -72 29 -71 33
rect -67 29 -65 33
rect -72 28 -65 29
rect -63 31 -55 34
rect 6 38 13 39
rect 6 34 7 38
rect 11 34 13 38
rect 6 33 13 34
rect -63 28 -53 31
rect -61 22 -53 28
rect -51 22 -46 31
rect -44 30 -37 31
rect 8 30 13 33
rect 15 34 20 39
rect 90 38 97 39
rect 90 34 91 38
rect 95 34 97 38
rect 15 30 29 34
rect -44 26 -42 30
rect -38 26 -37 30
rect -44 25 -37 26
rect 20 26 21 30
rect 25 26 29 30
rect 20 25 29 26
rect 31 33 39 34
rect 31 29 33 33
rect 37 29 39 33
rect 31 25 39 29
rect 41 31 49 34
rect 41 27 43 31
rect 47 27 49 31
rect 41 25 49 27
rect -44 22 -39 25
rect -61 21 -55 22
rect -61 17 -60 21
rect -56 17 -55 21
rect -61 16 -55 17
rect 44 22 49 25
rect 51 22 56 34
rect 58 22 66 34
rect 90 33 97 34
rect 92 30 97 33
rect 99 34 104 39
rect 99 30 113 34
rect 104 26 105 30
rect 109 26 113 30
rect 104 25 113 26
rect 115 33 123 34
rect 115 29 117 33
rect 121 29 123 33
rect 115 25 123 29
rect 125 31 133 34
rect 125 27 127 31
rect 131 27 133 31
rect 125 25 133 27
rect 60 21 66 22
rect 60 17 61 21
rect 65 17 66 21
rect 60 16 66 17
rect 128 22 133 25
rect 135 22 140 34
rect 142 22 150 34
rect 160 33 167 34
rect 160 29 161 33
rect 165 29 167 33
rect 160 28 167 29
rect 169 31 177 34
rect 169 28 179 31
rect 171 22 179 28
rect 181 22 186 31
rect 188 30 195 31
rect 188 26 190 30
rect 194 26 195 30
rect 188 25 195 26
rect 188 22 193 25
rect 144 21 150 22
rect 144 17 145 21
rect 149 17 150 21
rect 144 16 150 17
rect 171 21 177 22
rect 171 17 172 21
rect 176 17 177 21
rect 171 16 177 17
rect 21 -1 28 0
rect 21 -5 22 -1
rect 26 -5 28 -1
rect 21 -6 28 -5
rect 30 -1 38 0
rect 30 -5 32 -1
rect 36 -5 38 -1
rect 30 -6 38 -5
rect 40 -1 48 0
rect 40 -5 42 -1
rect 46 -5 48 -1
rect 40 -6 48 -5
rect 50 -1 57 0
rect 50 -5 52 -1
rect 56 -5 57 -1
rect 50 -6 57 -5
<< pdiffusion >>
rect -70 57 -65 63
rect -72 56 -65 57
rect -72 52 -71 56
rect -67 52 -65 56
rect -72 51 -65 52
rect -63 61 -57 63
rect -63 56 -55 61
rect -63 52 -61 56
rect -57 52 -55 56
rect -63 51 -55 52
rect -53 56 -45 61
rect -53 52 -51 56
rect -47 52 -45 56
rect -53 51 -45 52
rect -43 60 -36 61
rect -43 56 -41 60
rect -37 56 -36 60
rect 16 58 21 79
rect -43 51 -36 56
rect 14 57 21 58
rect 14 53 15 57
rect 19 53 21 57
rect 14 52 21 53
rect 23 78 35 79
rect 23 74 25 78
rect 29 74 35 78
rect 23 71 35 74
rect 23 67 25 71
rect 29 70 35 71
rect 52 70 57 79
rect 29 67 37 70
rect 23 52 37 67
rect 39 57 47 70
rect 39 53 41 57
rect 45 53 47 57
rect 39 52 47 53
rect 49 64 57 70
rect 49 60 51 64
rect 55 60 57 64
rect 49 52 57 60
rect 59 73 64 79
rect 59 72 66 73
rect 59 68 61 72
rect 65 68 66 72
rect 59 67 66 68
rect 59 52 64 67
rect 100 58 105 79
rect 98 57 105 58
rect 98 53 99 57
rect 103 53 105 57
rect 98 52 105 53
rect 107 78 119 79
rect 107 74 109 78
rect 113 74 119 78
rect 107 71 119 74
rect 107 67 109 71
rect 113 70 119 71
rect 136 70 141 79
rect 113 67 121 70
rect 107 52 121 67
rect 123 57 131 70
rect 123 53 125 57
rect 129 53 131 57
rect 123 52 131 53
rect 133 64 141 70
rect 133 60 135 64
rect 139 60 141 64
rect 133 52 141 60
rect 143 73 148 79
rect 143 72 150 73
rect 143 68 145 72
rect 149 68 150 72
rect 143 67 150 68
rect 143 52 148 67
rect 162 57 167 63
rect 160 56 167 57
rect 160 52 161 56
rect 165 52 167 56
rect 160 51 167 52
rect 169 61 175 63
rect 169 56 177 61
rect 169 52 171 56
rect 175 52 177 56
rect 169 51 177 52
rect 179 56 187 61
rect 179 52 181 56
rect 185 52 187 56
rect 179 51 187 52
rect 189 60 196 61
rect 189 56 191 60
rect 195 56 196 60
rect 189 51 196 56
rect 40 -33 48 -30
rect 23 -38 28 -33
rect 21 -39 28 -38
rect 21 -43 22 -39
rect 26 -43 28 -39
rect 21 -44 28 -43
rect 23 -51 28 -44
rect 30 -51 35 -33
rect 37 -42 48 -33
rect 50 -36 55 -30
rect 50 -37 57 -36
rect 50 -41 52 -37
rect 56 -41 57 -37
rect 50 -42 57 -41
rect 37 -46 46 -42
rect 37 -50 40 -46
rect 44 -50 46 -46
rect 37 -51 46 -50
<< metal1 >>
rect -106 81 200 85
rect -106 77 -70 81
rect -66 77 -56 81
rect -52 77 -42 81
rect -38 78 41 81
rect -38 77 25 78
rect -106 -34 -102 77
rect -72 57 -68 64
rect -72 56 -67 57
rect -72 52 -71 56
rect -64 56 -60 77
rect -57 71 -44 72
rect -57 67 -54 71
rect -50 67 -48 71
rect -57 66 -44 67
rect -57 59 -51 66
rect -41 60 -37 77
rect 29 77 41 78
rect 45 78 125 81
rect 45 77 109 78
rect 6 66 18 72
rect 25 71 29 74
rect 113 77 125 78
rect 129 77 162 81
rect 166 77 176 81
rect 180 77 190 81
rect 194 77 200 81
rect 39 68 61 72
rect 65 68 66 72
rect 90 71 102 72
rect 39 67 43 68
rect 25 66 29 67
rect 6 63 11 66
rect 6 62 7 63
rect -64 52 -61 56
rect -57 52 -56 56
rect -52 52 -51 56
rect -47 52 -46 56
rect -41 55 -37 56
rect -2 59 7 62
rect 32 63 43 67
rect 90 67 95 71
rect 99 67 102 71
rect 90 66 102 67
rect 109 71 113 74
rect 123 68 145 72
rect 149 68 150 72
rect 123 67 127 68
rect 109 66 113 67
rect 32 59 36 63
rect 50 60 51 64
rect 55 60 66 64
rect -72 51 -67 52
rect -72 43 -68 51
rect -52 47 -46 52
rect -65 43 -64 47
rect -60 43 -46 47
rect -40 45 -36 48
rect -2 45 1 59
rect 6 58 11 59
rect 15 57 36 59
rect -72 34 -68 39
rect -72 33 -67 34
rect -72 29 -71 33
rect -67 29 -60 32
rect -72 26 -60 29
rect -56 30 -52 43
rect 7 53 15 54
rect 19 55 36 57
rect 7 50 19 53
rect -40 39 -36 41
rect -49 35 -45 39
rect -41 35 -36 39
rect -49 34 -36 35
rect 7 38 11 50
rect 32 48 36 55
rect 40 53 41 57
rect 45 56 46 57
rect 45 53 57 56
rect 40 52 57 53
rect 53 49 57 52
rect 53 48 58 49
rect 21 42 27 47
rect 32 44 44 48
rect 48 44 49 48
rect 53 44 54 48
rect 21 40 23 42
rect 14 38 23 40
rect 53 43 58 44
rect 62 44 66 60
rect 90 63 95 66
rect 90 59 91 63
rect 116 63 127 67
rect 116 59 120 63
rect 134 60 135 64
rect 139 60 150 64
rect 90 58 95 59
rect 99 57 120 59
rect 91 53 99 54
rect 103 55 120 57
rect 91 50 103 53
rect 53 39 57 43
rect 14 34 27 38
rect 33 35 57 39
rect 62 40 64 44
rect 7 33 11 34
rect 33 33 37 35
rect -56 26 -42 30
rect -38 26 -37 30
rect 20 26 21 30
rect 25 26 26 30
rect 62 31 66 40
rect 91 38 95 50
rect 116 48 120 55
rect 124 53 125 57
rect 129 56 130 57
rect 129 53 141 56
rect 124 52 141 53
rect 137 49 141 52
rect 137 48 142 49
rect 105 42 111 47
rect 116 44 128 48
rect 132 44 133 48
rect 137 44 138 48
rect 105 40 107 42
rect 98 38 107 40
rect 137 43 142 44
rect 137 39 141 43
rect 98 34 111 38
rect 117 35 141 39
rect 91 33 95 34
rect 117 33 121 35
rect 33 28 37 29
rect 42 27 43 31
rect 47 27 66 31
rect 20 21 26 26
rect 104 26 105 30
rect 109 26 110 30
rect 146 31 150 60
rect 160 57 164 64
rect 160 56 165 57
rect 160 52 161 56
rect 168 56 172 77
rect 175 71 188 72
rect 175 67 178 71
rect 182 67 184 71
rect 175 66 188 67
rect 175 59 181 66
rect 191 60 195 77
rect 168 52 171 56
rect 175 52 176 56
rect 180 52 181 56
rect 185 52 186 56
rect 191 55 195 56
rect 160 51 165 52
rect 160 43 164 51
rect 180 47 186 52
rect 167 43 168 47
rect 172 43 186 47
rect 192 46 196 48
rect 117 28 121 29
rect 126 27 127 31
rect 131 27 150 31
rect 154 40 164 43
rect 154 28 157 40
rect 104 21 110 26
rect 160 34 164 40
rect 160 33 165 34
rect 160 29 161 33
rect 165 29 172 32
rect 160 26 172 29
rect 176 30 180 43
rect 192 39 196 42
rect 183 35 187 39
rect 191 35 196 39
rect 183 34 196 35
rect 176 26 190 30
rect 194 26 195 30
rect -73 17 -70 21
rect -66 17 -60 21
rect -56 17 8 21
rect 12 17 61 21
rect 65 17 92 21
rect 96 17 145 21
rect 149 17 162 21
rect 166 17 172 21
rect 176 17 200 21
rect -73 13 200 17
rect 17 11 61 13
rect 17 7 23 11
rect 27 7 51 11
rect 55 7 61 11
rect 21 -1 27 7
rect 21 -5 22 -1
rect 26 -5 27 -1
rect 32 -1 36 0
rect 41 -1 47 7
rect 41 -5 42 -1
rect 46 -5 47 -1
rect 52 -1 57 2
rect 56 -5 57 -1
rect 32 -8 36 -5
rect 52 -6 57 -5
rect 32 -12 49 -8
rect 21 -24 25 -14
rect 29 -19 34 -15
rect 45 -16 49 -12
rect 29 -27 35 -23
rect 39 -27 42 -23
rect -107 -54 -102 -34
rect 29 -33 33 -27
rect 45 -31 49 -20
rect 16 -36 33 -33
rect 37 -35 49 -31
rect 37 -39 41 -35
rect 53 -36 57 -6
rect 52 -37 57 -36
rect 21 -43 22 -39
rect 26 -43 41 -39
rect 44 -41 52 -39
rect 56 -41 57 -37
rect 44 -43 57 -41
rect 39 -49 40 -46
rect 17 -50 40 -49
rect 44 -49 45 -46
rect 44 -50 51 -49
rect 17 -53 51 -50
rect 55 -53 61 -49
rect 17 -54 61 -53
rect -107 -57 61 -54
rect -107 -58 17 -57
<< metal2 >>
rect -44 68 21 71
rect -79 40 -72 43
rect -79 -25 -76 40
rect -36 41 -3 44
rect 17 44 20 68
rect 99 68 184 71
rect 68 40 101 43
rect 81 36 84 40
rect 193 36 196 42
rect 81 33 196 36
rect 157 24 158 27
rect 155 -24 158 24
rect -79 -28 15 -25
rect 25 -27 168 -24
rect 12 -32 15 -28
<< ntransistor >>
rect -65 28 -63 34
rect -53 22 -51 31
rect -46 22 -44 31
rect 13 30 15 39
rect 29 25 31 34
rect 39 25 41 34
rect 49 22 51 34
rect 56 22 58 34
rect 97 30 99 39
rect 113 25 115 34
rect 123 25 125 34
rect 133 22 135 34
rect 140 22 142 34
rect 167 28 169 34
rect 179 22 181 31
rect 186 22 188 31
rect 28 -6 30 0
rect 38 -6 40 0
rect 48 -6 50 0
<< ptransistor >>
rect -65 51 -63 63
rect -55 51 -53 61
rect -45 51 -43 61
rect 21 52 23 79
rect 37 52 39 70
rect 47 52 49 70
rect 57 52 59 79
rect 105 52 107 79
rect 121 52 123 70
rect 131 52 133 70
rect 141 52 143 79
rect 167 51 169 63
rect 177 51 179 61
rect 187 51 189 61
rect 28 -51 30 -33
rect 35 -51 37 -33
rect 48 -42 50 -30
<< polycontact >>
rect -54 67 -50 71
rect 7 59 11 63
rect -64 43 -60 47
rect 91 59 95 63
rect 44 44 48 48
rect 54 44 58 48
rect 178 67 182 71
rect -45 35 -41 39
rect 23 38 27 42
rect 128 44 132 48
rect 138 44 142 48
rect 168 43 172 47
rect 107 38 111 42
rect 187 35 191 39
rect 25 -19 29 -15
rect 37 -19 41 -15
rect 45 -20 49 -16
rect 35 -27 39 -23
<< ndcontact >>
rect -71 29 -67 33
rect 7 34 11 38
rect 91 34 95 38
rect -42 26 -38 30
rect 21 26 25 30
rect 33 29 37 33
rect 43 27 47 31
rect -60 17 -56 21
rect 105 26 109 30
rect 117 29 121 33
rect 127 27 131 31
rect 61 17 65 21
rect 161 29 165 33
rect 190 26 194 30
rect 145 17 149 21
rect 172 17 176 21
rect 22 -5 26 -1
rect 32 -5 36 -1
rect 42 -5 46 -1
rect 52 -5 56 -1
<< pdcontact >>
rect -71 52 -67 56
rect -61 52 -57 56
rect -51 52 -47 56
rect -41 56 -37 60
rect 15 53 19 57
rect 25 74 29 78
rect 25 67 29 71
rect 41 53 45 57
rect 51 60 55 64
rect 61 68 65 72
rect 99 53 103 57
rect 109 74 113 78
rect 109 67 113 71
rect 125 53 129 57
rect 135 60 139 64
rect 145 68 149 72
rect 161 52 165 56
rect 171 52 175 56
rect 181 52 185 56
rect 191 56 195 60
rect 22 -43 26 -39
rect 52 -41 56 -37
rect 40 -50 44 -46
<< m2contact >>
rect -48 67 -44 71
rect 95 67 99 71
rect -72 39 -68 43
rect -40 41 -36 45
rect -3 41 1 45
rect 17 40 21 44
rect 64 40 68 44
rect 101 40 105 44
rect 184 67 188 71
rect 153 24 157 28
rect 192 42 196 46
rect 21 -28 25 -24
rect 12 -36 16 -32
<< psubstratepcontact >>
rect -70 17 -66 21
rect 8 17 12 21
rect 92 17 96 21
rect 162 17 166 21
rect 23 7 27 11
rect 51 7 55 11
<< nsubstratencontact >>
rect -70 77 -66 81
rect -56 77 -52 81
rect -42 77 -38 81
rect 41 77 45 81
rect 125 77 129 81
rect 162 77 166 81
rect 176 77 180 81
rect 190 77 194 81
rect 51 -53 55 -49
<< psubstratepdiff >>
rect -71 21 -65 22
rect -71 17 -70 21
rect -66 17 -65 21
rect -71 16 -65 17
rect 7 21 13 22
rect 7 17 8 21
rect 12 17 13 21
rect 7 16 13 17
rect 91 21 97 22
rect 91 17 92 21
rect 96 17 97 21
rect 91 16 97 17
rect 161 21 167 22
rect 161 17 162 21
rect 166 17 167 21
rect 161 16 167 17
rect 22 11 56 12
rect 22 7 23 11
rect 27 7 51 11
rect 55 7 56 11
rect 22 6 56 7
<< nsubstratendiff >>
rect -71 81 -37 82
rect -71 77 -70 81
rect -66 77 -56 81
rect -52 77 -42 81
rect -38 77 -37 81
rect 40 81 46 82
rect -71 76 -37 77
rect 40 77 41 81
rect 45 77 46 81
rect 124 81 130 82
rect 40 76 46 77
rect 124 77 125 81
rect 129 77 130 81
rect 161 81 195 82
rect 124 76 130 77
rect 161 77 162 81
rect 166 77 176 81
rect 180 77 190 81
rect 194 77 195 81
rect 161 76 195 77
rect 50 -49 56 -48
rect 50 -53 51 -49
rect 55 -53 56 -49
rect 50 -54 56 -53
<< labels >>
rlabel polycontact 46 46 46 46 6 bn
rlabel ntransistor 57 33 57 33 6 an
rlabel metal1 16 37 16 37 6 a
rlabel metal1 9 43 9 43 6 bn
rlabel metal1 8 65 8 65 6 b
rlabel metal1 16 69 16 69 6 b
rlabel polycontact 24 41 24 41 6 a
rlabel metal1 36 17 36 17 6 vss
rlabel metal1 35 33 35 33 6 an
rlabel metal1 40 46 40 46 6 bn
rlabel metal1 36 81 36 81 6 vdd
rlabel polycontact 55 46 55 46 6 an
rlabel metal1 48 54 48 54 6 an
rlabel metal1 52 70 52 70 6 bn
rlabel metal1 120 17 120 17 6 vss
rlabel metal1 120 81 120 81 6 vdd
rlabel metal1 64 49 64 49 1 so
rlabel metal1 148 49 148 49 1 sum
rlabel ntransistor 141 33 141 33 1 son
rlabel metal1 136 70 136 70 1 cn
rlabel metal1 -54 17 -54 17 6 vss
rlabel metal1 -54 81 -54 81 6 vdd
rlabel metal1 178 81 178 81 6 vdd
rlabel metal1 178 17 178 17 6 vss
rlabel metal1 100 69 100 69 1 c
rlabel metal1 39 11 39 11 2 vss
rlabel metal1 39 -53 39 -53 2 vdd
rlabel metal1 -49 49 -49 49 1 co_n
rlabel metal1 -62 29 -62 29 1 co
rlabel metal1 162 45 162 45 1 c1
rlabel metal1 176 45 176 45 1 zc1_n
rlabel metal1 47 -21 47 -21 1 cout_n
rlabel metal1 55 -17 55 -17 1 cout
<< end >>
