magic
tech scmos
timestamp 1523022893
<< pwell >>
rect 2 379 20 383
rect 0 375 20 379
rect 0 339 48 375
rect 87 339 135 375
rect 180 339 228 375
rect 420 341 468 377
rect 513 341 561 377
rect 600 341 648 377
rect -71 216 72 252
rect 84 216 202 252
rect 258 218 401 254
rect 413 218 531 254
rect 585 221 728 257
rect 740 221 858 257
rect 15 190 63 216
rect 344 192 392 218
rect 671 195 719 221
rect -72 70 71 106
rect 83 70 201 106
rect 257 72 400 108
rect 412 72 530 108
rect 584 75 727 111
rect 739 75 857 111
rect 14 44 62 70
rect 343 46 391 72
rect 670 49 718 75
rect 215 -78 263 -42
rect 308 -78 356 -42
rect 395 -78 443 -42
<< nwell >>
rect 0 296 48 339
rect 87 296 135 339
rect 180 296 228 339
rect 420 304 468 341
rect 513 304 561 341
rect 420 301 561 304
rect 416 298 561 301
rect 600 310 648 341
rect 600 301 661 310
rect 600 298 728 301
rect -71 252 72 296
rect 84 295 228 296
rect 84 252 202 295
rect 258 254 401 298
rect 413 284 728 298
rect 413 254 531 284
rect 585 257 728 284
rect 740 257 858 301
rect 15 183 63 190
rect 344 185 392 192
rect 671 188 719 195
rect 11 170 63 183
rect 340 172 392 185
rect 667 175 719 188
rect 15 154 63 170
rect 344 156 392 172
rect 671 162 719 175
rect 4 150 70 154
rect 334 152 400 156
rect 642 155 753 162
rect -72 106 71 150
rect 83 106 201 150
rect 257 108 400 152
rect 412 108 530 152
rect 584 146 857 155
rect 584 111 727 146
rect 739 111 857 146
rect 14 37 62 44
rect 343 39 391 46
rect 670 42 718 49
rect 10 24 62 37
rect 339 26 391 39
rect 666 29 718 42
rect 14 0 62 24
rect 343 16 391 26
rect 217 2 449 16
rect 670 5 718 29
rect 215 -1 449 2
rect 215 -42 263 -1
rect 308 -42 356 -1
rect 395 -42 443 -1
<< polysilicon >>
rect 13 358 15 363
rect 20 358 22 363
rect 33 356 35 360
rect 100 358 102 363
rect 107 358 109 363
rect 120 356 122 360
rect 193 358 195 363
rect 200 358 202 363
rect 213 356 215 360
rect 433 358 435 362
rect 446 360 448 365
rect 453 360 455 365
rect 526 358 528 362
rect 539 360 541 365
rect 546 360 548 365
rect 613 358 615 362
rect 626 360 628 365
rect 633 360 635 365
rect 13 334 15 347
rect 20 342 22 347
rect 33 342 35 347
rect 19 341 25 342
rect 19 337 20 341
rect 24 337 25 341
rect 19 336 25 337
rect 29 341 35 342
rect 29 337 30 341
rect 34 337 35 341
rect 29 336 35 337
rect 9 333 15 334
rect 9 329 10 333
rect 14 329 15 333
rect 9 328 15 329
rect 13 325 15 328
rect 23 325 25 336
rect 33 332 35 336
rect 100 334 102 347
rect 107 342 109 347
rect 120 342 122 347
rect 106 341 112 342
rect 106 337 107 341
rect 111 337 112 341
rect 106 336 112 337
rect 116 341 122 342
rect 116 337 117 341
rect 121 337 122 341
rect 116 336 122 337
rect 96 333 102 334
rect 96 329 97 333
rect 101 329 102 333
rect 96 328 102 329
rect 100 325 102 328
rect 110 325 112 336
rect 120 332 122 336
rect 193 334 195 347
rect 200 342 202 347
rect 213 342 215 347
rect 199 341 205 342
rect 199 337 200 341
rect 204 337 205 341
rect 199 336 205 337
rect 209 341 215 342
rect 209 337 210 341
rect 214 337 215 341
rect 209 336 215 337
rect 189 333 195 334
rect 13 307 15 312
rect 23 307 25 312
rect 33 310 35 314
rect 189 329 190 333
rect 194 329 195 333
rect 189 328 195 329
rect 193 325 195 328
rect 203 325 205 336
rect 213 332 215 336
rect 433 344 435 349
rect 446 344 448 349
rect 433 343 439 344
rect 433 339 434 343
rect 438 339 439 343
rect 433 338 439 339
rect 443 343 449 344
rect 443 339 444 343
rect 448 339 449 343
rect 443 338 449 339
rect 433 334 435 338
rect 100 307 102 312
rect 110 307 112 312
rect 120 310 122 314
rect 443 327 445 338
rect 453 336 455 349
rect 526 344 528 349
rect 539 344 541 349
rect 526 343 532 344
rect 526 339 527 343
rect 531 339 532 343
rect 526 338 532 339
rect 536 343 542 344
rect 536 339 537 343
rect 541 339 542 343
rect 536 338 542 339
rect 453 335 459 336
rect 453 331 454 335
rect 458 331 459 335
rect 526 334 528 338
rect 453 330 459 331
rect 453 327 455 330
rect 193 307 195 312
rect 203 307 205 312
rect 213 310 215 314
rect 433 312 435 316
rect 536 327 538 338
rect 546 336 548 349
rect 613 344 615 349
rect 626 344 628 349
rect 613 343 619 344
rect 613 339 614 343
rect 618 339 619 343
rect 613 338 619 339
rect 623 343 629 344
rect 623 339 624 343
rect 628 339 629 343
rect 623 338 629 339
rect 546 335 552 336
rect 546 331 547 335
rect 551 331 552 335
rect 613 334 615 338
rect 546 330 552 331
rect 546 327 548 330
rect 443 309 445 314
rect 453 309 455 314
rect 526 312 528 316
rect 623 327 625 338
rect 633 336 635 349
rect 633 335 639 336
rect 633 331 634 335
rect 638 331 639 335
rect 633 330 639 331
rect 633 327 635 330
rect 536 309 538 314
rect 546 309 548 314
rect 613 312 615 316
rect 623 309 625 314
rect 633 309 635 314
rect 21 286 23 290
rect -55 278 -49 279
rect -65 270 -63 275
rect -55 274 -54 278
rect -50 274 -49 278
rect -55 273 -49 274
rect -55 268 -53 273
rect -45 268 -43 273
rect 6 270 12 271
rect 6 266 7 270
rect 11 266 12 270
rect 6 265 12 266
rect -65 255 -63 258
rect -55 255 -53 258
rect -65 254 -59 255
rect -65 250 -64 254
rect -60 250 -59 254
rect -55 252 -51 255
rect -65 249 -59 250
rect -65 241 -63 249
rect -53 238 -51 252
rect -45 247 -43 258
rect 10 256 12 265
rect 57 286 59 290
rect 105 286 107 290
rect 37 277 39 281
rect 47 277 49 281
rect 90 270 96 271
rect 90 266 91 270
rect 95 266 96 270
rect 90 265 96 266
rect 21 256 23 259
rect 37 256 39 259
rect 47 256 49 259
rect 57 256 59 259
rect 10 254 23 256
rect 29 254 39 256
rect 43 255 49 256
rect -46 246 -40 247
rect 13 246 15 254
rect 29 250 31 254
rect 43 251 44 255
rect 48 251 49 255
rect 43 250 49 251
rect 53 255 59 256
rect 53 251 54 255
rect 58 251 59 255
rect 94 256 96 265
rect 141 286 143 290
rect 121 277 123 281
rect 131 277 133 281
rect 350 288 352 292
rect 274 280 280 281
rect 177 278 183 279
rect 167 270 169 275
rect 177 274 178 278
rect 182 274 183 278
rect 177 273 183 274
rect 105 256 107 259
rect 121 256 123 259
rect 131 256 133 259
rect 141 256 143 259
rect 177 268 179 273
rect 187 268 189 273
rect 264 272 266 277
rect 274 276 275 280
rect 279 276 280 280
rect 274 275 280 276
rect 274 270 276 275
rect 284 270 286 275
rect 335 272 341 273
rect 335 268 336 272
rect 340 268 341 272
rect 335 267 341 268
rect 94 254 107 256
rect 113 254 123 256
rect 127 255 133 256
rect 53 250 59 251
rect 22 249 31 250
rect -46 242 -45 246
rect -41 242 -40 246
rect -46 241 -40 242
rect -46 238 -44 241
rect -65 231 -63 235
rect 22 245 23 249
rect 27 245 31 249
rect 47 246 49 250
rect 22 244 31 245
rect 29 241 31 244
rect 39 241 41 246
rect 47 244 51 246
rect 49 241 51 244
rect 56 241 58 250
rect 97 246 99 254
rect 113 250 115 254
rect 127 251 128 255
rect 132 251 133 255
rect 127 250 133 251
rect 137 255 143 256
rect 137 251 138 255
rect 142 251 143 255
rect 137 250 143 251
rect 167 255 169 258
rect 177 255 179 258
rect 167 254 173 255
rect 167 250 168 254
rect 172 250 173 254
rect 177 252 181 255
rect 106 249 115 250
rect 13 234 15 237
rect 13 232 18 234
rect -53 224 -51 229
rect -46 224 -44 229
rect 16 224 18 232
rect 29 228 31 232
rect 39 224 41 232
rect 106 245 107 249
rect 111 245 115 249
rect 131 246 133 250
rect 106 244 115 245
rect 113 241 115 244
rect 123 241 125 246
rect 131 244 135 246
rect 133 241 135 244
rect 140 241 142 250
rect 167 249 173 250
rect 167 241 169 249
rect 97 234 99 237
rect 97 232 102 234
rect 49 224 51 229
rect 56 224 58 229
rect 16 222 41 224
rect 100 224 102 232
rect 113 228 115 232
rect 123 224 125 232
rect 179 238 181 252
rect 187 247 189 258
rect 264 257 266 260
rect 274 257 276 260
rect 264 256 270 257
rect 264 252 265 256
rect 269 252 270 256
rect 274 254 278 257
rect 264 251 270 252
rect 186 246 192 247
rect 186 242 187 246
rect 191 242 192 246
rect 264 243 266 251
rect 186 241 192 242
rect 186 238 188 241
rect 167 231 169 235
rect 276 240 278 254
rect 284 249 286 260
rect 339 258 341 267
rect 386 288 388 292
rect 434 288 436 292
rect 366 279 368 283
rect 376 279 378 283
rect 419 272 425 273
rect 419 268 420 272
rect 424 268 425 272
rect 419 267 425 268
rect 350 258 352 261
rect 366 258 368 261
rect 376 258 378 261
rect 386 258 388 261
rect 339 256 352 258
rect 358 256 368 258
rect 372 257 378 258
rect 283 248 289 249
rect 342 248 344 256
rect 358 252 360 256
rect 372 253 373 257
rect 377 253 378 257
rect 372 252 378 253
rect 382 257 388 258
rect 382 253 383 257
rect 387 253 388 257
rect 423 258 425 267
rect 470 288 472 292
rect 450 279 452 283
rect 460 279 462 283
rect 677 291 679 295
rect 601 283 607 284
rect 506 280 512 281
rect 496 272 498 277
rect 506 276 507 280
rect 511 276 512 280
rect 506 275 512 276
rect 591 275 593 280
rect 601 279 602 283
rect 606 279 607 283
rect 601 278 607 279
rect 434 258 436 261
rect 450 258 452 261
rect 460 258 462 261
rect 470 258 472 261
rect 506 270 508 275
rect 516 270 518 275
rect 601 273 603 278
rect 611 273 613 278
rect 662 275 668 276
rect 662 271 663 275
rect 667 271 668 275
rect 662 270 668 271
rect 591 260 593 263
rect 601 260 603 263
rect 423 256 436 258
rect 442 256 452 258
rect 456 257 462 258
rect 382 252 388 253
rect 351 251 360 252
rect 283 244 284 248
rect 288 244 289 248
rect 283 243 289 244
rect 283 240 285 243
rect 264 233 266 237
rect 351 247 352 251
rect 356 247 360 251
rect 376 248 378 252
rect 351 246 360 247
rect 358 243 360 246
rect 368 243 370 248
rect 376 246 380 248
rect 378 243 380 246
rect 385 243 387 252
rect 426 248 428 256
rect 442 252 444 256
rect 456 253 457 257
rect 461 253 462 257
rect 456 252 462 253
rect 466 257 472 258
rect 466 253 467 257
rect 471 253 472 257
rect 466 252 472 253
rect 496 257 498 260
rect 506 257 508 260
rect 496 256 502 257
rect 496 252 497 256
rect 501 252 502 256
rect 506 254 510 257
rect 435 251 444 252
rect 342 236 344 239
rect 342 234 347 236
rect 133 224 135 229
rect 140 224 142 229
rect 100 222 125 224
rect 179 224 181 229
rect 186 224 188 229
rect 276 226 278 231
rect 283 226 285 231
rect 345 226 347 234
rect 358 230 360 234
rect 368 226 370 234
rect 435 247 436 251
rect 440 247 444 251
rect 460 248 462 252
rect 435 246 444 247
rect 442 243 444 246
rect 452 243 454 248
rect 460 246 464 248
rect 462 243 464 246
rect 469 243 471 252
rect 496 251 502 252
rect 496 243 498 251
rect 426 236 428 239
rect 426 234 431 236
rect 378 226 380 231
rect 385 226 387 231
rect 345 224 370 226
rect 429 226 431 234
rect 442 230 444 234
rect 452 226 454 234
rect 508 240 510 254
rect 516 249 518 260
rect 591 259 597 260
rect 591 255 592 259
rect 596 255 597 259
rect 601 257 605 260
rect 591 254 597 255
rect 515 248 521 249
rect 515 244 516 248
rect 520 244 521 248
rect 591 246 593 254
rect 515 243 521 244
rect 515 240 517 243
rect 603 243 605 257
rect 611 252 613 263
rect 666 261 668 270
rect 713 291 715 295
rect 761 291 763 295
rect 693 282 695 286
rect 703 282 705 286
rect 746 275 752 276
rect 746 271 747 275
rect 751 271 752 275
rect 746 270 752 271
rect 677 261 679 264
rect 693 261 695 264
rect 703 261 705 264
rect 713 261 715 264
rect 666 259 679 261
rect 685 259 695 261
rect 699 260 705 261
rect 610 251 616 252
rect 669 251 671 259
rect 685 255 687 259
rect 699 256 700 260
rect 704 256 705 260
rect 699 255 705 256
rect 709 260 715 261
rect 709 256 710 260
rect 714 256 715 260
rect 750 261 752 270
rect 797 291 799 295
rect 777 282 779 286
rect 787 282 789 286
rect 833 283 839 284
rect 823 275 825 280
rect 833 279 834 283
rect 838 279 839 283
rect 833 278 839 279
rect 761 261 763 264
rect 777 261 779 264
rect 787 261 789 264
rect 797 261 799 264
rect 833 273 835 278
rect 843 273 845 278
rect 750 259 763 261
rect 769 259 779 261
rect 783 260 789 261
rect 709 255 715 256
rect 678 254 687 255
rect 610 247 611 251
rect 615 247 616 251
rect 610 246 616 247
rect 610 243 612 246
rect 496 233 498 237
rect 591 236 593 240
rect 678 250 679 254
rect 683 250 687 254
rect 703 251 705 255
rect 678 249 687 250
rect 685 246 687 249
rect 695 246 697 251
rect 703 249 707 251
rect 705 246 707 249
rect 712 246 714 255
rect 753 251 755 259
rect 769 255 771 259
rect 783 256 784 260
rect 788 256 789 260
rect 783 255 789 256
rect 793 260 799 261
rect 793 256 794 260
rect 798 256 799 260
rect 793 255 799 256
rect 823 260 825 263
rect 833 260 835 263
rect 823 259 829 260
rect 823 255 824 259
rect 828 255 829 259
rect 833 257 837 260
rect 762 254 771 255
rect 669 239 671 242
rect 669 237 674 239
rect 462 226 464 231
rect 469 226 471 231
rect 429 224 454 226
rect 508 226 510 231
rect 515 226 517 231
rect 603 229 605 234
rect 610 229 612 234
rect 672 229 674 237
rect 685 233 687 237
rect 695 229 697 237
rect 762 250 763 254
rect 767 250 771 254
rect 787 251 789 255
rect 762 249 771 250
rect 769 246 771 249
rect 779 246 781 251
rect 787 249 791 251
rect 789 246 791 249
rect 796 246 798 255
rect 823 254 829 255
rect 823 246 825 254
rect 753 239 755 242
rect 753 237 758 239
rect 705 229 707 234
rect 712 229 714 234
rect 672 227 697 229
rect 756 229 758 237
rect 769 233 771 237
rect 779 229 781 237
rect 835 243 837 257
rect 843 252 845 263
rect 842 251 848 252
rect 842 247 843 251
rect 847 247 848 251
rect 842 246 848 247
rect 842 243 844 246
rect 823 236 825 240
rect 789 229 791 234
rect 796 229 798 234
rect 756 227 781 229
rect 835 229 837 234
rect 842 229 844 234
rect 28 207 30 211
rect 38 207 40 211
rect 48 207 50 211
rect 357 209 359 213
rect 367 209 369 213
rect 377 209 379 213
rect 684 212 686 216
rect 694 212 696 216
rect 704 212 706 216
rect 28 193 30 201
rect 24 192 30 193
rect 38 192 40 201
rect 48 192 50 201
rect 357 195 359 203
rect 24 188 25 192
rect 29 188 30 192
rect 44 191 50 192
rect 24 187 30 188
rect 28 174 30 187
rect 38 185 40 188
rect 44 187 45 191
rect 49 187 50 191
rect 353 194 359 195
rect 367 194 369 203
rect 377 194 379 203
rect 684 198 686 206
rect 353 190 354 194
rect 358 190 359 194
rect 373 193 379 194
rect 353 189 359 190
rect 44 186 50 187
rect 34 184 40 185
rect 34 180 35 184
rect 39 180 40 184
rect 34 179 40 180
rect 35 174 37 179
rect 48 177 50 186
rect 357 176 359 189
rect 367 187 369 190
rect 373 189 374 193
rect 378 189 379 193
rect 680 197 686 198
rect 694 197 696 206
rect 704 197 706 206
rect 680 193 681 197
rect 685 193 686 197
rect 700 196 706 197
rect 680 192 686 193
rect 373 188 379 189
rect 363 186 369 187
rect 363 182 364 186
rect 368 182 369 186
rect 363 181 369 182
rect 364 176 366 181
rect 377 179 379 188
rect 684 179 686 192
rect 694 190 696 193
rect 700 192 701 196
rect 705 192 706 196
rect 700 191 706 192
rect 690 189 696 190
rect 690 185 691 189
rect 695 185 696 189
rect 690 184 696 185
rect 691 179 693 184
rect 704 182 706 191
rect 48 161 50 165
rect 377 163 379 167
rect 704 166 706 170
rect 28 152 30 156
rect 35 152 37 156
rect 357 154 359 158
rect 364 154 366 158
rect 684 157 686 161
rect 691 157 693 161
rect 20 140 22 144
rect -56 132 -50 133
rect -66 124 -64 129
rect -56 128 -55 132
rect -51 128 -50 132
rect -56 127 -50 128
rect -56 122 -54 127
rect -46 122 -44 127
rect 5 124 11 125
rect 5 120 6 124
rect 10 120 11 124
rect 5 119 11 120
rect -66 109 -64 112
rect -56 109 -54 112
rect -66 108 -60 109
rect -66 104 -65 108
rect -61 104 -60 108
rect -56 106 -52 109
rect -66 103 -60 104
rect -66 95 -64 103
rect -54 92 -52 106
rect -46 101 -44 112
rect 9 110 11 119
rect 56 140 58 144
rect 104 140 106 144
rect 36 131 38 135
rect 46 131 48 135
rect 89 124 95 125
rect 89 120 90 124
rect 94 120 95 124
rect 89 119 95 120
rect 20 110 22 113
rect 36 110 38 113
rect 46 110 48 113
rect 56 110 58 113
rect 9 108 22 110
rect 28 108 38 110
rect 42 109 48 110
rect -47 100 -41 101
rect 12 100 14 108
rect 28 104 30 108
rect 42 105 43 109
rect 47 105 48 109
rect 42 104 48 105
rect 52 109 58 110
rect 52 105 53 109
rect 57 105 58 109
rect 93 110 95 119
rect 140 140 142 144
rect 120 131 122 135
rect 130 131 132 135
rect 349 142 351 146
rect 273 134 279 135
rect 176 132 182 133
rect 166 124 168 129
rect 176 128 177 132
rect 181 128 182 132
rect 176 127 182 128
rect 104 110 106 113
rect 120 110 122 113
rect 130 110 132 113
rect 140 110 142 113
rect 176 122 178 127
rect 186 122 188 127
rect 263 126 265 131
rect 273 130 274 134
rect 278 130 279 134
rect 273 129 279 130
rect 273 124 275 129
rect 283 124 285 129
rect 334 126 340 127
rect 334 122 335 126
rect 339 122 340 126
rect 334 121 340 122
rect 93 108 106 110
rect 112 108 122 110
rect 126 109 132 110
rect 52 104 58 105
rect 21 103 30 104
rect -47 96 -46 100
rect -42 96 -41 100
rect -47 95 -41 96
rect -47 92 -45 95
rect -66 85 -64 89
rect 21 99 22 103
rect 26 99 30 103
rect 46 100 48 104
rect 21 98 30 99
rect 28 95 30 98
rect 38 95 40 100
rect 46 98 50 100
rect 48 95 50 98
rect 55 95 57 104
rect 96 100 98 108
rect 112 104 114 108
rect 126 105 127 109
rect 131 105 132 109
rect 126 104 132 105
rect 136 109 142 110
rect 136 105 137 109
rect 141 105 142 109
rect 136 104 142 105
rect 166 109 168 112
rect 176 109 178 112
rect 166 108 172 109
rect 166 104 167 108
rect 171 104 172 108
rect 176 106 180 109
rect 105 103 114 104
rect 12 88 14 91
rect 12 86 17 88
rect -54 78 -52 83
rect -47 78 -45 83
rect 15 78 17 86
rect 28 82 30 86
rect 38 78 40 86
rect 105 99 106 103
rect 110 99 114 103
rect 130 100 132 104
rect 105 98 114 99
rect 112 95 114 98
rect 122 95 124 100
rect 130 98 134 100
rect 132 95 134 98
rect 139 95 141 104
rect 166 103 172 104
rect 166 95 168 103
rect 96 88 98 91
rect 96 86 101 88
rect 48 78 50 83
rect 55 78 57 83
rect 15 76 40 78
rect 99 78 101 86
rect 112 82 114 86
rect 122 78 124 86
rect 178 92 180 106
rect 186 101 188 112
rect 263 111 265 114
rect 273 111 275 114
rect 263 110 269 111
rect 263 106 264 110
rect 268 106 269 110
rect 273 108 277 111
rect 263 105 269 106
rect 185 100 191 101
rect 185 96 186 100
rect 190 96 191 100
rect 263 97 265 105
rect 185 95 191 96
rect 185 92 187 95
rect 166 85 168 89
rect 275 94 277 108
rect 283 103 285 114
rect 338 112 340 121
rect 385 142 387 146
rect 433 142 435 146
rect 365 133 367 137
rect 375 133 377 137
rect 418 126 424 127
rect 418 122 419 126
rect 423 122 424 126
rect 418 121 424 122
rect 349 112 351 115
rect 365 112 367 115
rect 375 112 377 115
rect 385 112 387 115
rect 338 110 351 112
rect 357 110 367 112
rect 371 111 377 112
rect 282 102 288 103
rect 341 102 343 110
rect 357 106 359 110
rect 371 107 372 111
rect 376 107 377 111
rect 371 106 377 107
rect 381 111 387 112
rect 381 107 382 111
rect 386 107 387 111
rect 422 112 424 121
rect 469 142 471 146
rect 449 133 451 137
rect 459 133 461 137
rect 676 145 678 149
rect 600 137 606 138
rect 505 134 511 135
rect 495 126 497 131
rect 505 130 506 134
rect 510 130 511 134
rect 505 129 511 130
rect 590 129 592 134
rect 600 133 601 137
rect 605 133 606 137
rect 600 132 606 133
rect 433 112 435 115
rect 449 112 451 115
rect 459 112 461 115
rect 469 112 471 115
rect 505 124 507 129
rect 515 124 517 129
rect 600 127 602 132
rect 610 127 612 132
rect 661 129 667 130
rect 661 125 662 129
rect 666 125 667 129
rect 661 124 667 125
rect 590 114 592 117
rect 600 114 602 117
rect 422 110 435 112
rect 441 110 451 112
rect 455 111 461 112
rect 381 106 387 107
rect 350 105 359 106
rect 282 98 283 102
rect 287 98 288 102
rect 282 97 288 98
rect 282 94 284 97
rect 263 87 265 91
rect 350 101 351 105
rect 355 101 359 105
rect 375 102 377 106
rect 350 100 359 101
rect 357 97 359 100
rect 367 97 369 102
rect 375 100 379 102
rect 377 97 379 100
rect 384 97 386 106
rect 425 102 427 110
rect 441 106 443 110
rect 455 107 456 111
rect 460 107 461 111
rect 455 106 461 107
rect 465 111 471 112
rect 465 107 466 111
rect 470 107 471 111
rect 465 106 471 107
rect 495 111 497 114
rect 505 111 507 114
rect 495 110 501 111
rect 495 106 496 110
rect 500 106 501 110
rect 505 108 509 111
rect 434 105 443 106
rect 341 90 343 93
rect 341 88 346 90
rect 132 78 134 83
rect 139 78 141 83
rect 99 76 124 78
rect 178 78 180 83
rect 185 78 187 83
rect 275 80 277 85
rect 282 80 284 85
rect 344 80 346 88
rect 357 84 359 88
rect 367 80 369 88
rect 434 101 435 105
rect 439 101 443 105
rect 459 102 461 106
rect 434 100 443 101
rect 441 97 443 100
rect 451 97 453 102
rect 459 100 463 102
rect 461 97 463 100
rect 468 97 470 106
rect 495 105 501 106
rect 495 97 497 105
rect 425 90 427 93
rect 425 88 430 90
rect 377 80 379 85
rect 384 80 386 85
rect 344 78 369 80
rect 428 80 430 88
rect 441 84 443 88
rect 451 80 453 88
rect 507 94 509 108
rect 515 103 517 114
rect 590 113 596 114
rect 590 109 591 113
rect 595 109 596 113
rect 600 111 604 114
rect 590 108 596 109
rect 514 102 520 103
rect 514 98 515 102
rect 519 98 520 102
rect 590 100 592 108
rect 514 97 520 98
rect 514 94 516 97
rect 602 97 604 111
rect 610 106 612 117
rect 665 115 667 124
rect 712 145 714 149
rect 760 145 762 149
rect 692 136 694 140
rect 702 136 704 140
rect 745 129 751 130
rect 745 125 746 129
rect 750 125 751 129
rect 745 124 751 125
rect 676 115 678 118
rect 692 115 694 118
rect 702 115 704 118
rect 712 115 714 118
rect 665 113 678 115
rect 684 113 694 115
rect 698 114 704 115
rect 609 105 615 106
rect 668 105 670 113
rect 684 109 686 113
rect 698 110 699 114
rect 703 110 704 114
rect 698 109 704 110
rect 708 114 714 115
rect 708 110 709 114
rect 713 110 714 114
rect 749 115 751 124
rect 796 145 798 149
rect 776 136 778 140
rect 786 136 788 140
rect 832 137 838 138
rect 822 129 824 134
rect 832 133 833 137
rect 837 133 838 137
rect 832 132 838 133
rect 760 115 762 118
rect 776 115 778 118
rect 786 115 788 118
rect 796 115 798 118
rect 832 127 834 132
rect 842 127 844 132
rect 749 113 762 115
rect 768 113 778 115
rect 782 114 788 115
rect 708 109 714 110
rect 677 108 686 109
rect 609 101 610 105
rect 614 101 615 105
rect 609 100 615 101
rect 609 97 611 100
rect 495 87 497 91
rect 590 90 592 94
rect 677 104 678 108
rect 682 104 686 108
rect 702 105 704 109
rect 677 103 686 104
rect 684 100 686 103
rect 694 100 696 105
rect 702 103 706 105
rect 704 100 706 103
rect 711 100 713 109
rect 752 105 754 113
rect 768 109 770 113
rect 782 110 783 114
rect 787 110 788 114
rect 782 109 788 110
rect 792 114 798 115
rect 792 110 793 114
rect 797 110 798 114
rect 792 109 798 110
rect 822 114 824 117
rect 832 114 834 117
rect 822 113 828 114
rect 822 109 823 113
rect 827 109 828 113
rect 832 111 836 114
rect 761 108 770 109
rect 668 93 670 96
rect 668 91 673 93
rect 461 80 463 85
rect 468 80 470 85
rect 428 78 453 80
rect 507 80 509 85
rect 514 80 516 85
rect 602 83 604 88
rect 609 83 611 88
rect 671 83 673 91
rect 684 87 686 91
rect 694 83 696 91
rect 761 104 762 108
rect 766 104 770 108
rect 786 105 788 109
rect 761 103 770 104
rect 768 100 770 103
rect 778 100 780 105
rect 786 103 790 105
rect 788 100 790 103
rect 795 100 797 109
rect 822 108 828 109
rect 822 100 824 108
rect 752 93 754 96
rect 752 91 757 93
rect 704 83 706 88
rect 711 83 713 88
rect 671 81 696 83
rect 755 83 757 91
rect 768 87 770 91
rect 778 83 780 91
rect 834 97 836 111
rect 842 106 844 117
rect 841 105 847 106
rect 841 101 842 105
rect 846 101 847 105
rect 841 100 847 101
rect 841 97 843 100
rect 822 90 824 94
rect 788 83 790 88
rect 795 83 797 88
rect 755 81 780 83
rect 834 83 836 88
rect 841 83 843 88
rect 27 61 29 65
rect 37 61 39 65
rect 47 61 49 65
rect 356 63 358 67
rect 366 63 368 67
rect 376 63 378 67
rect 683 66 685 70
rect 693 66 695 70
rect 703 66 705 70
rect 27 47 29 55
rect 23 46 29 47
rect 37 46 39 55
rect 47 46 49 55
rect 356 49 358 57
rect 23 42 24 46
rect 28 42 29 46
rect 43 45 49 46
rect 23 41 29 42
rect 27 28 29 41
rect 37 39 39 42
rect 43 41 44 45
rect 48 41 49 45
rect 352 48 358 49
rect 366 48 368 57
rect 376 48 378 57
rect 683 52 685 60
rect 352 44 353 48
rect 357 44 358 48
rect 372 47 378 48
rect 352 43 358 44
rect 43 40 49 41
rect 33 38 39 39
rect 33 34 34 38
rect 38 34 39 38
rect 33 33 39 34
rect 34 28 36 33
rect 47 31 49 40
rect 356 30 358 43
rect 366 41 368 44
rect 372 43 373 47
rect 377 43 378 47
rect 679 51 685 52
rect 693 51 695 60
rect 703 51 705 60
rect 679 47 680 51
rect 684 47 685 51
rect 699 50 705 51
rect 679 46 685 47
rect 372 42 378 43
rect 362 40 368 41
rect 362 36 363 40
rect 367 36 368 40
rect 362 35 368 36
rect 363 30 365 35
rect 376 33 378 42
rect 683 33 685 46
rect 693 44 695 47
rect 699 46 700 50
rect 704 46 705 50
rect 699 45 705 46
rect 689 43 695 44
rect 689 39 690 43
rect 694 39 695 43
rect 689 38 695 39
rect 690 33 692 38
rect 703 36 705 45
rect 47 15 49 19
rect 376 17 378 21
rect 703 20 705 24
rect 27 6 29 10
rect 34 6 36 10
rect 356 8 358 12
rect 363 8 365 12
rect 683 11 685 15
rect 690 11 692 15
rect 228 -17 230 -13
rect 238 -15 240 -10
rect 248 -15 250 -10
rect 321 -17 323 -13
rect 331 -15 333 -10
rect 341 -15 343 -10
rect 228 -39 230 -35
rect 238 -39 240 -28
rect 248 -31 250 -28
rect 248 -32 254 -31
rect 248 -36 249 -32
rect 253 -36 254 -32
rect 408 -17 410 -13
rect 418 -15 420 -10
rect 428 -15 430 -10
rect 248 -37 254 -36
rect 228 -40 234 -39
rect 228 -44 229 -40
rect 233 -44 234 -40
rect 228 -45 234 -44
rect 238 -40 244 -39
rect 238 -44 239 -40
rect 243 -44 244 -40
rect 238 -45 244 -44
rect 228 -50 230 -45
rect 241 -50 243 -45
rect 248 -50 250 -37
rect 321 -39 323 -35
rect 331 -39 333 -28
rect 341 -31 343 -28
rect 341 -32 347 -31
rect 341 -36 342 -32
rect 346 -36 347 -32
rect 341 -37 347 -36
rect 321 -40 327 -39
rect 321 -44 322 -40
rect 326 -44 327 -40
rect 321 -45 327 -44
rect 331 -40 337 -39
rect 331 -44 332 -40
rect 336 -44 337 -40
rect 331 -45 337 -44
rect 321 -50 323 -45
rect 334 -50 336 -45
rect 341 -50 343 -37
rect 408 -39 410 -35
rect 418 -39 420 -28
rect 428 -31 430 -28
rect 428 -32 434 -31
rect 428 -36 429 -32
rect 433 -36 434 -32
rect 428 -37 434 -36
rect 408 -40 414 -39
rect 408 -44 409 -40
rect 413 -44 414 -40
rect 408 -45 414 -44
rect 418 -40 424 -39
rect 418 -44 419 -40
rect 423 -44 424 -40
rect 418 -45 424 -44
rect 408 -50 410 -45
rect 421 -50 423 -45
rect 428 -50 430 -37
rect 228 -63 230 -59
rect 241 -66 243 -61
rect 248 -66 250 -61
rect 321 -63 323 -59
rect 334 -66 336 -61
rect 341 -66 343 -61
rect 408 -63 410 -59
rect 421 -66 423 -61
rect 428 -66 430 -61
<< ndiffusion >>
rect 24 367 31 368
rect 24 363 26 367
rect 30 363 31 367
rect 24 358 31 363
rect 111 367 118 368
rect 111 363 113 367
rect 117 363 118 367
rect 6 357 13 358
rect 6 353 7 357
rect 11 353 13 357
rect 6 352 13 353
rect 8 347 13 352
rect 15 347 20 358
rect 22 356 31 358
rect 111 358 118 363
rect 204 367 211 368
rect 204 363 206 367
rect 210 363 211 367
rect 93 357 100 358
rect 22 347 33 356
rect 35 355 42 356
rect 35 351 37 355
rect 41 351 42 355
rect 93 353 94 357
rect 98 353 100 357
rect 93 352 100 353
rect 35 350 42 351
rect 35 347 40 350
rect 95 347 100 352
rect 102 347 107 358
rect 109 356 118 358
rect 204 358 211 363
rect 437 369 444 370
rect 437 365 438 369
rect 442 365 444 369
rect 186 357 193 358
rect 109 347 120 356
rect 122 355 129 356
rect 122 351 124 355
rect 128 351 129 355
rect 186 353 187 357
rect 191 353 193 357
rect 186 352 193 353
rect 122 350 129 351
rect 122 347 127 350
rect 188 347 193 352
rect 195 347 200 358
rect 202 356 211 358
rect 437 360 444 365
rect 530 369 537 370
rect 530 365 531 369
rect 535 365 537 369
rect 437 358 446 360
rect 426 357 433 358
rect 202 347 213 356
rect 215 355 222 356
rect 215 351 217 355
rect 221 351 222 355
rect 426 353 427 357
rect 431 353 433 357
rect 426 352 433 353
rect 215 350 222 351
rect 215 347 220 350
rect 428 349 433 352
rect 435 349 446 358
rect 448 349 453 360
rect 455 359 462 360
rect 455 355 457 359
rect 461 355 462 359
rect 530 360 537 365
rect 617 369 624 370
rect 617 365 618 369
rect 622 365 624 369
rect 530 358 539 360
rect 455 354 462 355
rect 519 357 526 358
rect 455 349 460 354
rect 519 353 520 357
rect 524 353 526 357
rect 519 352 526 353
rect 521 349 526 352
rect 528 349 539 358
rect 541 349 546 360
rect 548 359 555 360
rect 548 355 550 359
rect 554 355 555 359
rect 617 360 624 365
rect 617 358 626 360
rect 548 354 555 355
rect 606 357 613 358
rect 548 349 553 354
rect 606 353 607 357
rect 611 353 613 357
rect 606 352 613 353
rect 608 349 613 352
rect 615 349 626 358
rect 628 349 633 360
rect 635 359 642 360
rect 635 355 637 359
rect 641 355 642 359
rect 635 354 642 355
rect 635 349 640 354
rect -72 240 -65 241
rect -72 236 -71 240
rect -67 236 -65 240
rect -72 235 -65 236
rect -63 238 -55 241
rect 6 245 13 246
rect 6 241 7 245
rect 11 241 13 245
rect 6 240 13 241
rect -63 235 -53 238
rect -61 229 -53 235
rect -51 229 -46 238
rect -44 237 -37 238
rect 8 237 13 240
rect 15 241 20 246
rect 90 245 97 246
rect 90 241 91 245
rect 95 241 97 245
rect 15 237 29 241
rect -44 233 -42 237
rect -38 233 -37 237
rect -44 232 -37 233
rect 20 233 21 237
rect 25 233 29 237
rect 20 232 29 233
rect 31 240 39 241
rect 31 236 33 240
rect 37 236 39 240
rect 31 232 39 236
rect 41 238 49 241
rect 41 234 43 238
rect 47 234 49 238
rect 41 232 49 234
rect -44 229 -39 232
rect -61 228 -55 229
rect -61 224 -60 228
rect -56 224 -55 228
rect -61 223 -55 224
rect 44 229 49 232
rect 51 229 56 241
rect 58 229 66 241
rect 90 240 97 241
rect 92 237 97 240
rect 99 241 104 246
rect 99 237 113 241
rect 104 233 105 237
rect 109 233 113 237
rect 104 232 113 233
rect 115 240 123 241
rect 115 236 117 240
rect 121 236 123 240
rect 115 232 123 236
rect 125 238 133 241
rect 125 234 127 238
rect 131 234 133 238
rect 125 232 133 234
rect 60 228 66 229
rect 60 224 61 228
rect 65 224 66 228
rect 60 223 66 224
rect 128 229 133 232
rect 135 229 140 241
rect 142 229 150 241
rect 160 240 167 241
rect 160 236 161 240
rect 165 236 167 240
rect 160 235 167 236
rect 169 238 177 241
rect 257 242 264 243
rect 257 238 258 242
rect 262 238 264 242
rect 169 235 179 238
rect 171 229 179 235
rect 181 229 186 238
rect 188 237 195 238
rect 257 237 264 238
rect 266 240 274 243
rect 335 247 342 248
rect 335 243 336 247
rect 340 243 342 247
rect 335 242 342 243
rect 266 237 276 240
rect 188 233 190 237
rect 194 233 195 237
rect 188 232 195 233
rect 188 229 193 232
rect 268 231 276 237
rect 278 231 283 240
rect 285 239 292 240
rect 337 239 342 242
rect 344 243 349 248
rect 419 247 426 248
rect 419 243 420 247
rect 424 243 426 247
rect 344 239 358 243
rect 285 235 287 239
rect 291 235 292 239
rect 285 234 292 235
rect 349 235 350 239
rect 354 235 358 239
rect 349 234 358 235
rect 360 242 368 243
rect 360 238 362 242
rect 366 238 368 242
rect 360 234 368 238
rect 370 240 378 243
rect 370 236 372 240
rect 376 236 378 240
rect 370 234 378 236
rect 285 231 290 234
rect 144 228 150 229
rect 144 224 145 228
rect 149 224 150 228
rect 144 223 150 224
rect 171 228 177 229
rect 171 224 172 228
rect 176 224 177 228
rect 268 230 274 231
rect 268 226 269 230
rect 273 226 274 230
rect 268 225 274 226
rect 373 231 378 234
rect 380 231 385 243
rect 387 231 395 243
rect 419 242 426 243
rect 421 239 426 242
rect 428 243 433 248
rect 428 239 442 243
rect 433 235 434 239
rect 438 235 442 239
rect 433 234 442 235
rect 444 242 452 243
rect 444 238 446 242
rect 450 238 452 242
rect 444 234 452 238
rect 454 240 462 243
rect 454 236 456 240
rect 460 236 462 240
rect 454 234 462 236
rect 389 230 395 231
rect 389 226 390 230
rect 394 226 395 230
rect 389 225 395 226
rect 457 231 462 234
rect 464 231 469 243
rect 471 231 479 243
rect 489 242 496 243
rect 489 238 490 242
rect 494 238 496 242
rect 489 237 496 238
rect 498 240 506 243
rect 584 245 591 246
rect 584 241 585 245
rect 589 241 591 245
rect 584 240 591 241
rect 593 243 601 246
rect 662 250 669 251
rect 662 246 663 250
rect 667 246 669 250
rect 662 245 669 246
rect 593 240 603 243
rect 498 237 508 240
rect 500 231 508 237
rect 510 231 515 240
rect 517 239 524 240
rect 517 235 519 239
rect 523 235 524 239
rect 517 234 524 235
rect 595 234 603 240
rect 605 234 610 243
rect 612 242 619 243
rect 664 242 669 245
rect 671 246 676 251
rect 746 250 753 251
rect 746 246 747 250
rect 751 246 753 250
rect 671 242 685 246
rect 612 238 614 242
rect 618 238 619 242
rect 612 237 619 238
rect 676 238 677 242
rect 681 238 685 242
rect 676 237 685 238
rect 687 245 695 246
rect 687 241 689 245
rect 693 241 695 245
rect 687 237 695 241
rect 697 243 705 246
rect 697 239 699 243
rect 703 239 705 243
rect 697 237 705 239
rect 612 234 617 237
rect 517 231 522 234
rect 473 230 479 231
rect 473 226 474 230
rect 478 226 479 230
rect 473 225 479 226
rect 500 230 506 231
rect 500 226 501 230
rect 505 226 506 230
rect 595 233 601 234
rect 595 229 596 233
rect 600 229 601 233
rect 595 228 601 229
rect 700 234 705 237
rect 707 234 712 246
rect 714 234 722 246
rect 746 245 753 246
rect 748 242 753 245
rect 755 246 760 251
rect 755 242 769 246
rect 760 238 761 242
rect 765 238 769 242
rect 760 237 769 238
rect 771 245 779 246
rect 771 241 773 245
rect 777 241 779 245
rect 771 237 779 241
rect 781 243 789 246
rect 781 239 783 243
rect 787 239 789 243
rect 781 237 789 239
rect 716 233 722 234
rect 716 229 717 233
rect 721 229 722 233
rect 716 228 722 229
rect 784 234 789 237
rect 791 234 796 246
rect 798 234 806 246
rect 816 245 823 246
rect 816 241 817 245
rect 821 241 823 245
rect 816 240 823 241
rect 825 243 833 246
rect 825 240 835 243
rect 827 234 835 240
rect 837 234 842 243
rect 844 242 851 243
rect 844 238 846 242
rect 850 238 851 242
rect 844 237 851 238
rect 844 234 849 237
rect 800 233 806 234
rect 800 229 801 233
rect 805 229 806 233
rect 800 228 806 229
rect 827 233 833 234
rect 827 229 828 233
rect 832 229 833 233
rect 827 228 833 229
rect 500 225 506 226
rect 171 223 177 224
rect 677 211 684 212
rect 350 208 357 209
rect 21 206 28 207
rect 21 202 22 206
rect 26 202 28 206
rect 21 201 28 202
rect 30 206 38 207
rect 30 202 32 206
rect 36 202 38 206
rect 30 201 38 202
rect 40 206 48 207
rect 40 202 42 206
rect 46 202 48 206
rect 40 201 48 202
rect 50 206 57 207
rect 50 202 52 206
rect 56 202 57 206
rect 350 204 351 208
rect 355 204 357 208
rect 350 203 357 204
rect 359 208 367 209
rect 359 204 361 208
rect 365 204 367 208
rect 359 203 367 204
rect 369 208 377 209
rect 369 204 371 208
rect 375 204 377 208
rect 369 203 377 204
rect 379 208 386 209
rect 379 204 381 208
rect 385 204 386 208
rect 677 207 678 211
rect 682 207 684 211
rect 677 206 684 207
rect 686 211 694 212
rect 686 207 688 211
rect 692 207 694 211
rect 686 206 694 207
rect 696 211 704 212
rect 696 207 698 211
rect 702 207 704 211
rect 696 206 704 207
rect 706 211 713 212
rect 706 207 708 211
rect 712 207 713 211
rect 706 206 713 207
rect 379 203 386 204
rect 50 201 57 202
rect -73 94 -66 95
rect -73 90 -72 94
rect -68 90 -66 94
rect -73 89 -66 90
rect -64 92 -56 95
rect 5 99 12 100
rect 5 95 6 99
rect 10 95 12 99
rect 5 94 12 95
rect -64 89 -54 92
rect -62 83 -54 89
rect -52 83 -47 92
rect -45 91 -38 92
rect 7 91 12 94
rect 14 95 19 100
rect 89 99 96 100
rect 89 95 90 99
rect 94 95 96 99
rect 14 91 28 95
rect -45 87 -43 91
rect -39 87 -38 91
rect -45 86 -38 87
rect 19 87 20 91
rect 24 87 28 91
rect 19 86 28 87
rect 30 94 38 95
rect 30 90 32 94
rect 36 90 38 94
rect 30 86 38 90
rect 40 92 48 95
rect 40 88 42 92
rect 46 88 48 92
rect 40 86 48 88
rect -45 83 -40 86
rect -62 82 -56 83
rect -62 78 -61 82
rect -57 78 -56 82
rect -62 77 -56 78
rect 43 83 48 86
rect 50 83 55 95
rect 57 83 65 95
rect 89 94 96 95
rect 91 91 96 94
rect 98 95 103 100
rect 98 91 112 95
rect 103 87 104 91
rect 108 87 112 91
rect 103 86 112 87
rect 114 94 122 95
rect 114 90 116 94
rect 120 90 122 94
rect 114 86 122 90
rect 124 92 132 95
rect 124 88 126 92
rect 130 88 132 92
rect 124 86 132 88
rect 59 82 65 83
rect 59 78 60 82
rect 64 78 65 82
rect 59 77 65 78
rect 127 83 132 86
rect 134 83 139 95
rect 141 83 149 95
rect 159 94 166 95
rect 159 90 160 94
rect 164 90 166 94
rect 159 89 166 90
rect 168 92 176 95
rect 256 96 263 97
rect 256 92 257 96
rect 261 92 263 96
rect 168 89 178 92
rect 170 83 178 89
rect 180 83 185 92
rect 187 91 194 92
rect 256 91 263 92
rect 265 94 273 97
rect 334 101 341 102
rect 334 97 335 101
rect 339 97 341 101
rect 334 96 341 97
rect 265 91 275 94
rect 187 87 189 91
rect 193 87 194 91
rect 187 86 194 87
rect 187 83 192 86
rect 267 85 275 91
rect 277 85 282 94
rect 284 93 291 94
rect 336 93 341 96
rect 343 97 348 102
rect 418 101 425 102
rect 418 97 419 101
rect 423 97 425 101
rect 343 93 357 97
rect 284 89 286 93
rect 290 89 291 93
rect 284 88 291 89
rect 348 89 349 93
rect 353 89 357 93
rect 348 88 357 89
rect 359 96 367 97
rect 359 92 361 96
rect 365 92 367 96
rect 359 88 367 92
rect 369 94 377 97
rect 369 90 371 94
rect 375 90 377 94
rect 369 88 377 90
rect 284 85 289 88
rect 143 82 149 83
rect 143 78 144 82
rect 148 78 149 82
rect 143 77 149 78
rect 170 82 176 83
rect 170 78 171 82
rect 175 78 176 82
rect 267 84 273 85
rect 267 80 268 84
rect 272 80 273 84
rect 267 79 273 80
rect 372 85 377 88
rect 379 85 384 97
rect 386 85 394 97
rect 418 96 425 97
rect 420 93 425 96
rect 427 97 432 102
rect 427 93 441 97
rect 432 89 433 93
rect 437 89 441 93
rect 432 88 441 89
rect 443 96 451 97
rect 443 92 445 96
rect 449 92 451 96
rect 443 88 451 92
rect 453 94 461 97
rect 453 90 455 94
rect 459 90 461 94
rect 453 88 461 90
rect 388 84 394 85
rect 388 80 389 84
rect 393 80 394 84
rect 388 79 394 80
rect 456 85 461 88
rect 463 85 468 97
rect 470 85 478 97
rect 488 96 495 97
rect 488 92 489 96
rect 493 92 495 96
rect 488 91 495 92
rect 497 94 505 97
rect 583 99 590 100
rect 583 95 584 99
rect 588 95 590 99
rect 583 94 590 95
rect 592 97 600 100
rect 661 104 668 105
rect 661 100 662 104
rect 666 100 668 104
rect 661 99 668 100
rect 592 94 602 97
rect 497 91 507 94
rect 499 85 507 91
rect 509 85 514 94
rect 516 93 523 94
rect 516 89 518 93
rect 522 89 523 93
rect 516 88 523 89
rect 594 88 602 94
rect 604 88 609 97
rect 611 96 618 97
rect 663 96 668 99
rect 670 100 675 105
rect 745 104 752 105
rect 745 100 746 104
rect 750 100 752 104
rect 670 96 684 100
rect 611 92 613 96
rect 617 92 618 96
rect 611 91 618 92
rect 675 92 676 96
rect 680 92 684 96
rect 675 91 684 92
rect 686 99 694 100
rect 686 95 688 99
rect 692 95 694 99
rect 686 91 694 95
rect 696 97 704 100
rect 696 93 698 97
rect 702 93 704 97
rect 696 91 704 93
rect 611 88 616 91
rect 516 85 521 88
rect 472 84 478 85
rect 472 80 473 84
rect 477 80 478 84
rect 472 79 478 80
rect 499 84 505 85
rect 499 80 500 84
rect 504 80 505 84
rect 594 87 600 88
rect 594 83 595 87
rect 599 83 600 87
rect 594 82 600 83
rect 699 88 704 91
rect 706 88 711 100
rect 713 88 721 100
rect 745 99 752 100
rect 747 96 752 99
rect 754 100 759 105
rect 754 96 768 100
rect 759 92 760 96
rect 764 92 768 96
rect 759 91 768 92
rect 770 99 778 100
rect 770 95 772 99
rect 776 95 778 99
rect 770 91 778 95
rect 780 97 788 100
rect 780 93 782 97
rect 786 93 788 97
rect 780 91 788 93
rect 715 87 721 88
rect 715 83 716 87
rect 720 83 721 87
rect 715 82 721 83
rect 783 88 788 91
rect 790 88 795 100
rect 797 88 805 100
rect 815 99 822 100
rect 815 95 816 99
rect 820 95 822 99
rect 815 94 822 95
rect 824 97 832 100
rect 824 94 834 97
rect 826 88 834 94
rect 836 88 841 97
rect 843 96 850 97
rect 843 92 845 96
rect 849 92 850 96
rect 843 91 850 92
rect 843 88 848 91
rect 799 87 805 88
rect 799 83 800 87
rect 804 83 805 87
rect 799 82 805 83
rect 826 87 832 88
rect 826 83 827 87
rect 831 83 832 87
rect 826 82 832 83
rect 499 79 505 80
rect 170 77 176 78
rect 676 65 683 66
rect 349 62 356 63
rect 20 60 27 61
rect 20 56 21 60
rect 25 56 27 60
rect 20 55 27 56
rect 29 60 37 61
rect 29 56 31 60
rect 35 56 37 60
rect 29 55 37 56
rect 39 60 47 61
rect 39 56 41 60
rect 45 56 47 60
rect 39 55 47 56
rect 49 60 56 61
rect 49 56 51 60
rect 55 56 56 60
rect 349 58 350 62
rect 354 58 356 62
rect 349 57 356 58
rect 358 62 366 63
rect 358 58 360 62
rect 364 58 366 62
rect 358 57 366 58
rect 368 62 376 63
rect 368 58 370 62
rect 374 58 376 62
rect 368 57 376 58
rect 378 62 385 63
rect 378 58 380 62
rect 384 58 385 62
rect 676 61 677 65
rect 681 61 683 65
rect 676 60 683 61
rect 685 65 693 66
rect 685 61 687 65
rect 691 61 693 65
rect 685 60 693 61
rect 695 65 703 66
rect 695 61 697 65
rect 701 61 703 65
rect 695 60 703 61
rect 705 65 712 66
rect 705 61 707 65
rect 711 61 712 65
rect 705 60 712 61
rect 378 57 385 58
rect 49 55 56 56
rect 223 -53 228 -50
rect 221 -54 228 -53
rect 221 -58 222 -54
rect 226 -58 228 -54
rect 221 -59 228 -58
rect 230 -59 241 -50
rect 232 -61 241 -59
rect 243 -61 248 -50
rect 250 -55 255 -50
rect 316 -53 321 -50
rect 314 -54 321 -53
rect 250 -56 257 -55
rect 250 -60 252 -56
rect 256 -60 257 -56
rect 314 -58 315 -54
rect 319 -58 321 -54
rect 314 -59 321 -58
rect 323 -59 334 -50
rect 250 -61 257 -60
rect 232 -66 239 -61
rect 325 -61 334 -59
rect 336 -61 341 -50
rect 343 -55 348 -50
rect 403 -53 408 -50
rect 401 -54 408 -53
rect 343 -56 350 -55
rect 343 -60 345 -56
rect 349 -60 350 -56
rect 401 -58 402 -54
rect 406 -58 408 -54
rect 401 -59 408 -58
rect 410 -59 421 -50
rect 343 -61 350 -60
rect 232 -70 233 -66
rect 237 -70 239 -66
rect 232 -71 239 -70
rect 325 -66 332 -61
rect 412 -61 421 -59
rect 423 -61 428 -50
rect 430 -55 435 -50
rect 430 -56 437 -55
rect 430 -60 432 -56
rect 436 -60 437 -56
rect 430 -61 437 -60
rect 325 -70 326 -66
rect 330 -70 332 -66
rect 325 -71 332 -70
rect 412 -66 419 -61
rect 412 -70 413 -66
rect 417 -70 419 -66
rect 412 -71 419 -70
<< pdiffusion >>
rect 27 325 33 332
rect 6 317 13 325
rect 6 313 7 317
rect 11 313 13 317
rect 6 312 13 313
rect 15 324 23 325
rect 15 320 17 324
rect 21 320 23 324
rect 15 317 23 320
rect 15 313 17 317
rect 21 313 23 317
rect 15 312 23 313
rect 25 319 33 325
rect 25 315 27 319
rect 31 315 33 319
rect 25 314 33 315
rect 35 331 42 332
rect 35 327 37 331
rect 41 327 42 331
rect 35 324 42 327
rect 114 325 120 332
rect 35 320 37 324
rect 41 320 42 324
rect 35 319 42 320
rect 35 314 40 319
rect 93 317 100 325
rect 25 312 31 314
rect 93 313 94 317
rect 98 313 100 317
rect 93 312 100 313
rect 102 324 110 325
rect 102 320 104 324
rect 108 320 110 324
rect 102 317 110 320
rect 102 313 104 317
rect 108 313 110 317
rect 102 312 110 313
rect 112 319 120 325
rect 112 315 114 319
rect 118 315 120 319
rect 112 314 120 315
rect 122 331 129 332
rect 122 327 124 331
rect 128 327 129 331
rect 122 324 129 327
rect 426 333 433 334
rect 207 325 213 332
rect 122 320 124 324
rect 128 320 129 324
rect 122 319 129 320
rect 122 314 127 319
rect 186 317 193 325
rect 112 312 118 314
rect 186 313 187 317
rect 191 313 193 317
rect 186 312 193 313
rect 195 324 203 325
rect 195 320 197 324
rect 201 320 203 324
rect 195 317 203 320
rect 195 313 197 317
rect 201 313 203 317
rect 195 312 203 313
rect 205 319 213 325
rect 205 315 207 319
rect 211 315 213 319
rect 205 314 213 315
rect 215 331 222 332
rect 215 327 217 331
rect 221 327 222 331
rect 215 324 222 327
rect 215 320 217 324
rect 221 320 222 324
rect 426 329 427 333
rect 431 329 433 333
rect 426 326 433 329
rect 426 322 427 326
rect 431 322 433 326
rect 426 321 433 322
rect 215 319 222 320
rect 215 314 220 319
rect 428 316 433 321
rect 435 327 441 334
rect 519 333 526 334
rect 519 329 520 333
rect 524 329 526 333
rect 435 321 443 327
rect 435 317 437 321
rect 441 317 443 321
rect 435 316 443 317
rect 205 312 211 314
rect 437 314 443 316
rect 445 326 453 327
rect 445 322 447 326
rect 451 322 453 326
rect 445 319 453 322
rect 445 315 447 319
rect 451 315 453 319
rect 445 314 453 315
rect 455 319 462 327
rect 519 326 526 329
rect 519 322 520 326
rect 524 322 526 326
rect 519 321 526 322
rect 455 315 457 319
rect 461 315 462 319
rect 521 316 526 321
rect 528 327 534 334
rect 606 333 613 334
rect 606 329 607 333
rect 611 329 613 333
rect 528 321 536 327
rect 528 317 530 321
rect 534 317 536 321
rect 528 316 536 317
rect 455 314 462 315
rect 530 314 536 316
rect 538 326 546 327
rect 538 322 540 326
rect 544 322 546 326
rect 538 319 546 322
rect 538 315 540 319
rect 544 315 546 319
rect 538 314 546 315
rect 548 319 555 327
rect 606 326 613 329
rect 606 322 607 326
rect 611 322 613 326
rect 606 321 613 322
rect 548 315 550 319
rect 554 315 555 319
rect 608 316 613 321
rect 615 327 621 334
rect 615 321 623 327
rect 615 317 617 321
rect 621 317 623 321
rect 615 316 623 317
rect 548 314 555 315
rect 617 314 623 316
rect 625 326 633 327
rect 625 322 627 326
rect 631 322 633 326
rect 625 319 633 322
rect 625 315 627 319
rect 631 315 633 319
rect 625 314 633 315
rect 635 319 642 327
rect 635 315 637 319
rect 641 315 642 319
rect 635 314 642 315
rect -70 264 -65 270
rect -72 263 -65 264
rect -72 259 -71 263
rect -67 259 -65 263
rect -72 258 -65 259
rect -63 268 -57 270
rect -63 263 -55 268
rect -63 259 -61 263
rect -57 259 -55 263
rect -63 258 -55 259
rect -53 263 -45 268
rect -53 259 -51 263
rect -47 259 -45 263
rect -53 258 -45 259
rect -43 267 -36 268
rect -43 263 -41 267
rect -37 263 -36 267
rect 16 265 21 286
rect -43 258 -36 263
rect 14 264 21 265
rect 14 260 15 264
rect 19 260 21 264
rect 14 259 21 260
rect 23 285 35 286
rect 23 281 25 285
rect 29 281 35 285
rect 23 278 35 281
rect 23 274 25 278
rect 29 277 35 278
rect 52 277 57 286
rect 29 274 37 277
rect 23 259 37 274
rect 39 264 47 277
rect 39 260 41 264
rect 45 260 47 264
rect 39 259 47 260
rect 49 271 57 277
rect 49 267 51 271
rect 55 267 57 271
rect 49 259 57 267
rect 59 280 64 286
rect 59 279 66 280
rect 59 275 61 279
rect 65 275 66 279
rect 59 274 66 275
rect 59 259 64 274
rect 100 265 105 286
rect 98 264 105 265
rect 98 260 99 264
rect 103 260 105 264
rect 98 259 105 260
rect 107 285 119 286
rect 107 281 109 285
rect 113 281 119 285
rect 107 278 119 281
rect 107 274 109 278
rect 113 277 119 278
rect 136 277 141 286
rect 113 274 121 277
rect 107 259 121 274
rect 123 264 131 277
rect 123 260 125 264
rect 129 260 131 264
rect 123 259 131 260
rect 133 271 141 277
rect 133 267 135 271
rect 139 267 141 271
rect 133 259 141 267
rect 143 280 148 286
rect 143 279 150 280
rect 143 275 145 279
rect 149 275 150 279
rect 143 274 150 275
rect 143 259 148 274
rect 162 264 167 270
rect 160 263 167 264
rect 160 259 161 263
rect 165 259 167 263
rect 160 258 167 259
rect 169 268 175 270
rect 169 263 177 268
rect 169 259 171 263
rect 175 259 177 263
rect 169 258 177 259
rect 179 263 187 268
rect 179 259 181 263
rect 185 259 187 263
rect 179 258 187 259
rect 189 267 196 268
rect 189 263 191 267
rect 195 263 196 267
rect 259 266 264 272
rect 189 258 196 263
rect 257 265 264 266
rect 257 261 258 265
rect 262 261 264 265
rect 257 260 264 261
rect 266 270 272 272
rect 266 265 274 270
rect 266 261 268 265
rect 272 261 274 265
rect 266 260 274 261
rect 276 265 284 270
rect 276 261 278 265
rect 282 261 284 265
rect 276 260 284 261
rect 286 269 293 270
rect 286 265 288 269
rect 292 265 293 269
rect 345 267 350 288
rect 286 260 293 265
rect 343 266 350 267
rect 343 262 344 266
rect 348 262 350 266
rect 343 261 350 262
rect 352 287 364 288
rect 352 283 354 287
rect 358 283 364 287
rect 352 280 364 283
rect 352 276 354 280
rect 358 279 364 280
rect 381 279 386 288
rect 358 276 366 279
rect 352 261 366 276
rect 368 266 376 279
rect 368 262 370 266
rect 374 262 376 266
rect 368 261 376 262
rect 378 273 386 279
rect 378 269 380 273
rect 384 269 386 273
rect 378 261 386 269
rect 388 282 393 288
rect 388 281 395 282
rect 388 277 390 281
rect 394 277 395 281
rect 388 276 395 277
rect 388 261 393 276
rect 429 267 434 288
rect 427 266 434 267
rect 427 262 428 266
rect 432 262 434 266
rect 427 261 434 262
rect 436 287 448 288
rect 436 283 438 287
rect 442 283 448 287
rect 436 280 448 283
rect 436 276 438 280
rect 442 279 448 280
rect 465 279 470 288
rect 442 276 450 279
rect 436 261 450 276
rect 452 266 460 279
rect 452 262 454 266
rect 458 262 460 266
rect 452 261 460 262
rect 462 273 470 279
rect 462 269 464 273
rect 468 269 470 273
rect 462 261 470 269
rect 472 282 477 288
rect 472 281 479 282
rect 472 277 474 281
rect 478 277 479 281
rect 472 276 479 277
rect 472 261 477 276
rect 491 266 496 272
rect 489 265 496 266
rect 489 261 490 265
rect 494 261 496 265
rect 489 260 496 261
rect 498 270 504 272
rect 498 265 506 270
rect 498 261 500 265
rect 504 261 506 265
rect 498 260 506 261
rect 508 265 516 270
rect 508 261 510 265
rect 514 261 516 265
rect 508 260 516 261
rect 518 269 525 270
rect 586 269 591 275
rect 518 265 520 269
rect 524 265 525 269
rect 518 260 525 265
rect 584 268 591 269
rect 584 264 585 268
rect 589 264 591 268
rect 584 263 591 264
rect 593 273 599 275
rect 593 268 601 273
rect 593 264 595 268
rect 599 264 601 268
rect 593 263 601 264
rect 603 268 611 273
rect 603 264 605 268
rect 609 264 611 268
rect 603 263 611 264
rect 613 272 620 273
rect 613 268 615 272
rect 619 268 620 272
rect 672 270 677 291
rect 613 263 620 268
rect 670 269 677 270
rect 670 265 671 269
rect 675 265 677 269
rect 670 264 677 265
rect 679 290 691 291
rect 679 286 681 290
rect 685 286 691 290
rect 679 283 691 286
rect 679 279 681 283
rect 685 282 691 283
rect 708 282 713 291
rect 685 279 693 282
rect 679 264 693 279
rect 695 269 703 282
rect 695 265 697 269
rect 701 265 703 269
rect 695 264 703 265
rect 705 276 713 282
rect 705 272 707 276
rect 711 272 713 276
rect 705 264 713 272
rect 715 285 720 291
rect 715 284 722 285
rect 715 280 717 284
rect 721 280 722 284
rect 715 279 722 280
rect 715 264 720 279
rect 756 270 761 291
rect 754 269 761 270
rect 754 265 755 269
rect 759 265 761 269
rect 754 264 761 265
rect 763 290 775 291
rect 763 286 765 290
rect 769 286 775 290
rect 763 283 775 286
rect 763 279 765 283
rect 769 282 775 283
rect 792 282 797 291
rect 769 279 777 282
rect 763 264 777 279
rect 779 269 787 282
rect 779 265 781 269
rect 785 265 787 269
rect 779 264 787 265
rect 789 276 797 282
rect 789 272 791 276
rect 795 272 797 276
rect 789 264 797 272
rect 799 285 804 291
rect 799 284 806 285
rect 799 280 801 284
rect 805 280 806 284
rect 799 279 806 280
rect 799 264 804 279
rect 818 269 823 275
rect 816 268 823 269
rect 816 264 817 268
rect 821 264 823 268
rect 816 263 823 264
rect 825 273 831 275
rect 825 268 833 273
rect 825 264 827 268
rect 831 264 833 268
rect 825 263 833 264
rect 835 268 843 273
rect 835 264 837 268
rect 841 264 843 268
rect 835 263 843 264
rect 845 272 852 273
rect 845 268 847 272
rect 851 268 852 272
rect 845 263 852 268
rect 40 174 48 177
rect 23 169 28 174
rect 21 168 28 169
rect 21 164 22 168
rect 26 164 28 168
rect 21 163 28 164
rect 23 156 28 163
rect 30 156 35 174
rect 37 165 48 174
rect 50 171 55 177
rect 696 179 704 182
rect 369 176 377 179
rect 352 171 357 176
rect 50 170 57 171
rect 50 166 52 170
rect 56 166 57 170
rect 50 165 57 166
rect 350 170 357 171
rect 350 166 351 170
rect 355 166 357 170
rect 350 165 357 166
rect 37 161 46 165
rect 37 157 40 161
rect 44 157 46 161
rect 37 156 46 157
rect 352 158 357 165
rect 359 158 364 176
rect 366 167 377 176
rect 379 173 384 179
rect 679 174 684 179
rect 677 173 684 174
rect 379 172 386 173
rect 379 168 381 172
rect 385 168 386 172
rect 677 169 678 173
rect 682 169 684 173
rect 677 168 684 169
rect 379 167 386 168
rect 366 163 375 167
rect 366 159 369 163
rect 373 159 375 163
rect 679 161 684 168
rect 686 161 691 179
rect 693 170 704 179
rect 706 176 711 182
rect 706 175 713 176
rect 706 171 708 175
rect 712 171 713 175
rect 706 170 713 171
rect 693 166 702 170
rect 693 162 696 166
rect 700 162 702 166
rect 693 161 702 162
rect 366 158 375 159
rect -71 118 -66 124
rect -73 117 -66 118
rect -73 113 -72 117
rect -68 113 -66 117
rect -73 112 -66 113
rect -64 122 -58 124
rect -64 117 -56 122
rect -64 113 -62 117
rect -58 113 -56 117
rect -64 112 -56 113
rect -54 117 -46 122
rect -54 113 -52 117
rect -48 113 -46 117
rect -54 112 -46 113
rect -44 121 -37 122
rect -44 117 -42 121
rect -38 117 -37 121
rect 15 119 20 140
rect -44 112 -37 117
rect 13 118 20 119
rect 13 114 14 118
rect 18 114 20 118
rect 13 113 20 114
rect 22 139 34 140
rect 22 135 24 139
rect 28 135 34 139
rect 22 132 34 135
rect 22 128 24 132
rect 28 131 34 132
rect 51 131 56 140
rect 28 128 36 131
rect 22 113 36 128
rect 38 118 46 131
rect 38 114 40 118
rect 44 114 46 118
rect 38 113 46 114
rect 48 125 56 131
rect 48 121 50 125
rect 54 121 56 125
rect 48 113 56 121
rect 58 134 63 140
rect 58 133 65 134
rect 58 129 60 133
rect 64 129 65 133
rect 58 128 65 129
rect 58 113 63 128
rect 99 119 104 140
rect 97 118 104 119
rect 97 114 98 118
rect 102 114 104 118
rect 97 113 104 114
rect 106 139 118 140
rect 106 135 108 139
rect 112 135 118 139
rect 106 132 118 135
rect 106 128 108 132
rect 112 131 118 132
rect 135 131 140 140
rect 112 128 120 131
rect 106 113 120 128
rect 122 118 130 131
rect 122 114 124 118
rect 128 114 130 118
rect 122 113 130 114
rect 132 125 140 131
rect 132 121 134 125
rect 138 121 140 125
rect 132 113 140 121
rect 142 134 147 140
rect 142 133 149 134
rect 142 129 144 133
rect 148 129 149 133
rect 142 128 149 129
rect 142 113 147 128
rect 161 118 166 124
rect 159 117 166 118
rect 159 113 160 117
rect 164 113 166 117
rect 159 112 166 113
rect 168 122 174 124
rect 168 117 176 122
rect 168 113 170 117
rect 174 113 176 117
rect 168 112 176 113
rect 178 117 186 122
rect 178 113 180 117
rect 184 113 186 117
rect 178 112 186 113
rect 188 121 195 122
rect 188 117 190 121
rect 194 117 195 121
rect 258 120 263 126
rect 188 112 195 117
rect 256 119 263 120
rect 256 115 257 119
rect 261 115 263 119
rect 256 114 263 115
rect 265 124 271 126
rect 265 119 273 124
rect 265 115 267 119
rect 271 115 273 119
rect 265 114 273 115
rect 275 119 283 124
rect 275 115 277 119
rect 281 115 283 119
rect 275 114 283 115
rect 285 123 292 124
rect 285 119 287 123
rect 291 119 292 123
rect 344 121 349 142
rect 285 114 292 119
rect 342 120 349 121
rect 342 116 343 120
rect 347 116 349 120
rect 342 115 349 116
rect 351 141 363 142
rect 351 137 353 141
rect 357 137 363 141
rect 351 134 363 137
rect 351 130 353 134
rect 357 133 363 134
rect 380 133 385 142
rect 357 130 365 133
rect 351 115 365 130
rect 367 120 375 133
rect 367 116 369 120
rect 373 116 375 120
rect 367 115 375 116
rect 377 127 385 133
rect 377 123 379 127
rect 383 123 385 127
rect 377 115 385 123
rect 387 136 392 142
rect 387 135 394 136
rect 387 131 389 135
rect 393 131 394 135
rect 387 130 394 131
rect 387 115 392 130
rect 428 121 433 142
rect 426 120 433 121
rect 426 116 427 120
rect 431 116 433 120
rect 426 115 433 116
rect 435 141 447 142
rect 435 137 437 141
rect 441 137 447 141
rect 435 134 447 137
rect 435 130 437 134
rect 441 133 447 134
rect 464 133 469 142
rect 441 130 449 133
rect 435 115 449 130
rect 451 120 459 133
rect 451 116 453 120
rect 457 116 459 120
rect 451 115 459 116
rect 461 127 469 133
rect 461 123 463 127
rect 467 123 469 127
rect 461 115 469 123
rect 471 136 476 142
rect 471 135 478 136
rect 471 131 473 135
rect 477 131 478 135
rect 471 130 478 131
rect 471 115 476 130
rect 490 120 495 126
rect 488 119 495 120
rect 488 115 489 119
rect 493 115 495 119
rect 488 114 495 115
rect 497 124 503 126
rect 497 119 505 124
rect 497 115 499 119
rect 503 115 505 119
rect 497 114 505 115
rect 507 119 515 124
rect 507 115 509 119
rect 513 115 515 119
rect 507 114 515 115
rect 517 123 524 124
rect 585 123 590 129
rect 517 119 519 123
rect 523 119 524 123
rect 517 114 524 119
rect 583 122 590 123
rect 583 118 584 122
rect 588 118 590 122
rect 583 117 590 118
rect 592 127 598 129
rect 592 122 600 127
rect 592 118 594 122
rect 598 118 600 122
rect 592 117 600 118
rect 602 122 610 127
rect 602 118 604 122
rect 608 118 610 122
rect 602 117 610 118
rect 612 126 619 127
rect 612 122 614 126
rect 618 122 619 126
rect 671 124 676 145
rect 612 117 619 122
rect 669 123 676 124
rect 669 119 670 123
rect 674 119 676 123
rect 669 118 676 119
rect 678 144 690 145
rect 678 140 680 144
rect 684 140 690 144
rect 678 137 690 140
rect 678 133 680 137
rect 684 136 690 137
rect 707 136 712 145
rect 684 133 692 136
rect 678 118 692 133
rect 694 123 702 136
rect 694 119 696 123
rect 700 119 702 123
rect 694 118 702 119
rect 704 130 712 136
rect 704 126 706 130
rect 710 126 712 130
rect 704 118 712 126
rect 714 139 719 145
rect 714 138 721 139
rect 714 134 716 138
rect 720 134 721 138
rect 714 133 721 134
rect 714 118 719 133
rect 755 124 760 145
rect 753 123 760 124
rect 753 119 754 123
rect 758 119 760 123
rect 753 118 760 119
rect 762 144 774 145
rect 762 140 764 144
rect 768 140 774 144
rect 762 137 774 140
rect 762 133 764 137
rect 768 136 774 137
rect 791 136 796 145
rect 768 133 776 136
rect 762 118 776 133
rect 778 123 786 136
rect 778 119 780 123
rect 784 119 786 123
rect 778 118 786 119
rect 788 130 796 136
rect 788 126 790 130
rect 794 126 796 130
rect 788 118 796 126
rect 798 139 803 145
rect 798 138 805 139
rect 798 134 800 138
rect 804 134 805 138
rect 798 133 805 134
rect 798 118 803 133
rect 817 123 822 129
rect 815 122 822 123
rect 815 118 816 122
rect 820 118 822 122
rect 815 117 822 118
rect 824 127 830 129
rect 824 122 832 127
rect 824 118 826 122
rect 830 118 832 122
rect 824 117 832 118
rect 834 122 842 127
rect 834 118 836 122
rect 840 118 842 122
rect 834 117 842 118
rect 844 126 851 127
rect 844 122 846 126
rect 850 122 851 126
rect 844 117 851 122
rect 39 28 47 31
rect 22 23 27 28
rect 20 22 27 23
rect 20 18 21 22
rect 25 18 27 22
rect 20 17 27 18
rect 22 10 27 17
rect 29 10 34 28
rect 36 19 47 28
rect 49 25 54 31
rect 695 33 703 36
rect 368 30 376 33
rect 351 25 356 30
rect 49 24 56 25
rect 49 20 51 24
rect 55 20 56 24
rect 49 19 56 20
rect 349 24 356 25
rect 349 20 350 24
rect 354 20 356 24
rect 349 19 356 20
rect 36 15 45 19
rect 36 11 39 15
rect 43 11 45 15
rect 36 10 45 11
rect 351 12 356 19
rect 358 12 363 30
rect 365 21 376 30
rect 378 27 383 33
rect 678 28 683 33
rect 676 27 683 28
rect 378 26 385 27
rect 378 22 380 26
rect 384 22 385 26
rect 676 23 677 27
rect 681 23 683 27
rect 676 22 683 23
rect 378 21 385 22
rect 365 17 374 21
rect 365 13 368 17
rect 372 13 374 17
rect 678 15 683 22
rect 685 15 690 33
rect 692 24 703 33
rect 705 30 710 36
rect 705 29 712 30
rect 705 25 707 29
rect 711 25 712 29
rect 705 24 712 25
rect 692 20 701 24
rect 692 16 695 20
rect 699 16 701 20
rect 692 15 701 16
rect 365 12 374 13
rect 232 -17 238 -15
rect 223 -22 228 -17
rect 221 -23 228 -22
rect 221 -27 222 -23
rect 226 -27 228 -23
rect 221 -30 228 -27
rect 221 -34 222 -30
rect 226 -34 228 -30
rect 221 -35 228 -34
rect 230 -18 238 -17
rect 230 -22 232 -18
rect 236 -22 238 -18
rect 230 -28 238 -22
rect 240 -16 248 -15
rect 240 -20 242 -16
rect 246 -20 248 -16
rect 240 -23 248 -20
rect 240 -27 242 -23
rect 246 -27 248 -23
rect 240 -28 248 -27
rect 250 -16 257 -15
rect 250 -20 252 -16
rect 256 -20 257 -16
rect 325 -17 331 -15
rect 250 -28 257 -20
rect 316 -22 321 -17
rect 314 -23 321 -22
rect 314 -27 315 -23
rect 319 -27 321 -23
rect 230 -35 236 -28
rect 314 -30 321 -27
rect 314 -34 315 -30
rect 319 -34 321 -30
rect 314 -35 321 -34
rect 323 -18 331 -17
rect 323 -22 325 -18
rect 329 -22 331 -18
rect 323 -28 331 -22
rect 333 -16 341 -15
rect 333 -20 335 -16
rect 339 -20 341 -16
rect 333 -23 341 -20
rect 333 -27 335 -23
rect 339 -27 341 -23
rect 333 -28 341 -27
rect 343 -16 350 -15
rect 343 -20 345 -16
rect 349 -20 350 -16
rect 412 -17 418 -15
rect 343 -28 350 -20
rect 403 -22 408 -17
rect 401 -23 408 -22
rect 401 -27 402 -23
rect 406 -27 408 -23
rect 323 -35 329 -28
rect 401 -30 408 -27
rect 401 -34 402 -30
rect 406 -34 408 -30
rect 401 -35 408 -34
rect 410 -18 418 -17
rect 410 -22 412 -18
rect 416 -22 418 -18
rect 410 -28 418 -22
rect 420 -16 428 -15
rect 420 -20 422 -16
rect 426 -20 428 -16
rect 420 -23 428 -20
rect 420 -27 422 -23
rect 426 -27 428 -23
rect 420 -28 428 -27
rect 430 -16 437 -15
rect 430 -20 432 -16
rect 436 -20 437 -16
rect 430 -28 437 -20
rect 410 -35 416 -28
<< metal1 >>
rect -75 380 366 384
rect -75 358 -71 380
rect 7 371 8 374
rect 223 371 416 372
rect 422 371 466 373
rect 7 370 466 371
rect 515 370 559 373
rect 602 372 646 373
rect 602 370 654 372
rect 2 369 654 370
rect 2 367 428 369
rect 2 363 26 367
rect 30 363 36 367
rect 40 363 113 367
rect 117 363 123 367
rect 127 363 206 367
rect 210 363 216 367
rect 220 366 428 367
rect 220 363 226 366
rect 422 365 428 366
rect 432 365 438 369
rect 442 366 521 369
rect 442 365 466 366
rect 515 365 521 366
rect 525 365 531 369
rect 535 366 608 369
rect 535 365 559 366
rect 602 365 608 366
rect 612 365 618 369
rect 622 366 654 369
rect 622 365 646 366
rect 6 353 7 357
rect 11 353 26 357
rect -37 346 2 349
rect 6 346 18 350
rect -37 344 -34 346
rect -99 341 -34 344
rect 13 341 18 346
rect 22 349 26 353
rect 30 355 42 358
rect 30 352 37 355
rect 41 351 42 355
rect 93 353 94 357
rect 98 353 113 357
rect 37 350 42 351
rect 22 345 34 349
rect 30 341 34 345
rect 13 337 20 341
rect 24 337 27 341
rect 6 324 10 333
rect 14 329 19 333
rect 30 326 34 337
rect 38 336 42 350
rect 94 346 105 350
rect 100 341 105 346
rect 109 349 113 353
rect 117 355 129 358
rect 117 352 124 355
rect 128 351 129 355
rect 186 353 187 357
rect 191 353 206 357
rect 124 350 129 351
rect 109 345 121 349
rect 117 341 121 345
rect 100 337 107 341
rect 111 337 114 341
rect 38 333 67 336
rect 38 332 42 333
rect -1 320 10 324
rect 17 324 34 326
rect 21 322 34 324
rect 37 331 42 332
rect 41 327 42 331
rect 37 324 42 327
rect 17 317 21 320
rect 41 320 42 324
rect 37 319 42 320
rect 6 313 7 317
rect 11 313 12 317
rect 6 307 12 313
rect 17 312 21 313
rect 26 315 27 319
rect 31 315 32 319
rect 26 307 32 315
rect 2 303 36 307
rect 40 303 46 307
rect 2 299 46 303
rect 3 292 7 299
rect 63 297 67 333
rect 93 323 97 333
rect 101 329 106 333
rect 117 326 121 337
rect 125 332 129 350
rect 187 346 198 350
rect 193 341 198 346
rect 202 349 206 353
rect 210 355 222 358
rect 426 357 438 360
rect 210 352 217 355
rect 221 351 222 355
rect 235 351 304 355
rect 310 351 407 355
rect 412 351 413 355
rect 426 353 427 357
rect 431 354 438 357
rect 442 355 457 359
rect 461 355 462 359
rect 519 357 531 360
rect 426 352 431 353
rect 217 350 222 351
rect 202 345 214 349
rect 210 341 214 345
rect 193 337 200 341
rect 204 337 207 341
rect 90 320 97 323
rect 104 324 121 326
rect 108 322 121 324
rect 124 331 129 332
rect 128 327 129 331
rect 124 324 129 327
rect 104 317 108 320
rect 128 322 129 324
rect 128 320 135 322
rect 124 319 135 320
rect 186 323 190 333
rect 194 329 199 333
rect 210 326 214 337
rect 218 332 222 350
rect 426 345 430 352
rect 442 351 446 355
rect 519 353 520 357
rect 524 354 531 357
rect 535 355 550 359
rect 554 355 555 359
rect 606 357 618 360
rect 519 352 524 353
rect 370 341 430 345
rect 183 320 190 323
rect 197 324 214 326
rect 201 322 214 324
rect 217 331 222 332
rect 221 327 222 331
rect 235 329 292 332
rect 426 334 430 341
rect 434 347 446 351
rect 450 349 461 352
rect 434 343 438 347
rect 450 343 455 349
rect 441 339 444 343
rect 448 339 455 343
rect 519 341 523 352
rect 535 351 539 355
rect 606 353 607 357
rect 611 354 618 357
rect 622 355 637 359
rect 641 355 642 359
rect 606 352 611 353
rect 426 333 431 334
rect 298 329 408 332
rect 426 329 427 333
rect 217 324 222 327
rect 426 326 431 329
rect 93 313 94 317
rect 98 313 99 317
rect 93 307 99 313
rect 104 312 108 313
rect 113 315 114 319
rect 118 315 119 319
rect 197 317 201 320
rect 221 320 222 324
rect 217 319 222 320
rect 113 307 119 315
rect 186 313 187 317
rect 191 313 192 317
rect 186 307 192 313
rect 197 312 201 313
rect 206 315 207 319
rect 211 315 212 319
rect 426 322 427 326
rect 434 328 438 339
rect 496 338 523 341
rect 449 331 454 335
rect 434 326 451 328
rect 434 324 447 326
rect 426 321 431 322
rect 458 325 462 335
rect 496 326 500 338
rect 458 322 465 325
rect 206 307 212 315
rect 273 314 277 318
rect 436 317 437 321
rect 441 317 442 321
rect 235 311 409 314
rect 436 309 442 317
rect 447 319 451 322
rect 519 334 523 338
rect 527 347 539 351
rect 543 351 557 352
rect 543 349 554 351
rect 527 343 531 347
rect 543 343 548 349
rect 534 339 537 343
rect 541 339 548 343
rect 519 333 524 334
rect 519 329 520 333
rect 519 326 524 329
rect 519 322 520 326
rect 527 328 531 339
rect 606 338 610 352
rect 622 351 626 355
rect 542 331 547 335
rect 527 326 544 328
rect 527 324 540 326
rect 519 321 524 322
rect 551 325 555 335
rect 584 334 610 338
rect 614 347 626 351
rect 630 351 644 352
rect 630 349 641 351
rect 614 343 618 347
rect 630 343 635 349
rect 621 339 624 343
rect 628 339 635 343
rect 551 322 558 325
rect 570 324 571 328
rect 447 314 451 315
rect 456 315 457 319
rect 461 315 462 319
rect 456 309 462 315
rect 529 317 530 321
rect 534 317 535 321
rect 529 309 535 317
rect 540 319 544 322
rect 540 314 544 315
rect 549 315 550 319
rect 554 315 555 319
rect 549 309 555 315
rect 89 303 123 307
rect 127 303 133 307
rect 89 302 133 303
rect 182 303 216 307
rect 220 303 226 307
rect 89 299 116 302
rect 182 299 226 303
rect 422 305 428 309
rect 432 305 466 309
rect 515 305 521 309
rect 525 305 559 309
rect 422 301 466 305
rect 91 292 95 299
rect 128 295 161 298
rect 182 292 186 299
rect 458 297 462 301
rect 477 300 507 303
rect 515 301 559 305
rect 570 304 574 324
rect 416 296 520 297
rect 416 294 542 296
rect 551 294 555 301
rect 584 303 588 334
rect 606 333 611 334
rect 606 329 607 333
rect 594 304 598 324
rect 606 326 611 329
rect 606 322 607 326
rect 614 328 618 339
rect 629 331 634 335
rect 614 326 631 328
rect 614 324 627 326
rect 606 321 611 322
rect 638 326 642 335
rect 638 322 646 326
rect 616 317 617 321
rect 621 317 622 321
rect 616 309 622 317
rect 627 319 631 322
rect 627 314 631 315
rect 636 315 637 319
rect 641 315 642 319
rect 636 309 642 315
rect 602 305 608 309
rect 612 305 646 309
rect 602 301 646 305
rect 640 294 644 301
rect 654 294 856 297
rect 198 293 856 294
rect 198 292 586 293
rect -106 291 121 292
rect 134 291 586 292
rect -106 290 586 291
rect -106 288 259 290
rect -106 284 -70 288
rect -66 284 -56 288
rect -52 284 -42 288
rect -38 285 41 288
rect -38 284 25 285
rect -106 173 -102 284
rect -86 283 -71 284
rect -72 264 -68 271
rect -72 263 -67 264
rect -72 259 -71 263
rect -64 263 -60 284
rect -57 278 -44 279
rect -57 274 -54 278
rect -50 274 -48 278
rect -57 273 -44 274
rect -57 266 -51 273
rect -41 267 -37 284
rect 29 284 41 285
rect 45 285 125 288
rect 45 284 109 285
rect 6 273 18 279
rect 25 278 29 281
rect 113 284 125 285
rect 129 284 162 288
rect 166 284 176 288
rect 180 284 190 288
rect 194 286 259 288
rect 263 286 273 290
rect 277 286 287 290
rect 291 287 370 290
rect 291 286 354 287
rect 194 284 229 286
rect 39 275 61 279
rect 65 275 66 279
rect 90 278 102 279
rect 39 274 43 275
rect 25 273 29 274
rect 6 270 11 273
rect 6 269 7 270
rect -64 259 -61 263
rect -57 259 -56 263
rect -52 259 -51 263
rect -47 259 -46 263
rect -41 262 -37 263
rect -2 266 7 269
rect 32 270 43 274
rect 90 274 95 278
rect 99 274 102 278
rect 90 273 102 274
rect 109 278 113 281
rect 123 275 145 279
rect 149 275 150 279
rect 123 274 127 275
rect 109 273 113 274
rect 32 266 36 270
rect 50 267 51 271
rect 55 267 66 271
rect -72 258 -67 259
rect -72 250 -68 258
rect -52 254 -46 259
rect -65 250 -64 254
rect -60 250 -46 254
rect -40 252 -36 255
rect -2 252 1 266
rect 6 265 11 266
rect 15 264 36 266
rect -72 241 -68 246
rect -72 240 -67 241
rect -72 236 -71 240
rect -67 236 -60 239
rect -72 233 -60 236
rect -56 237 -52 250
rect 7 260 15 261
rect 19 262 36 264
rect 7 257 19 260
rect -40 246 -36 248
rect -49 242 -45 246
rect -41 242 -36 246
rect -49 241 -36 242
rect 7 245 11 257
rect 32 255 36 262
rect 40 260 41 264
rect 45 263 46 264
rect 45 260 57 263
rect 40 259 57 260
rect 53 256 57 259
rect 53 255 58 256
rect 21 249 27 254
rect 32 251 44 255
rect 48 251 49 255
rect 53 251 54 255
rect 21 247 23 249
rect 14 245 23 247
rect 53 250 58 251
rect 62 251 66 267
rect 90 270 95 273
rect 90 266 91 270
rect 116 270 127 274
rect 116 266 120 270
rect 134 267 135 271
rect 139 267 150 271
rect 90 265 95 266
rect 99 264 120 266
rect 91 260 99 261
rect 103 262 120 264
rect 91 257 103 260
rect 53 246 57 250
rect 14 241 27 245
rect 33 242 57 246
rect 62 247 64 251
rect 7 240 11 241
rect 33 240 37 242
rect -56 233 -42 237
rect -38 233 -37 237
rect 20 233 21 237
rect 25 233 26 237
rect 62 238 66 247
rect 91 245 95 257
rect 116 255 120 262
rect 124 260 125 264
rect 129 263 130 264
rect 129 260 141 263
rect 124 259 141 260
rect 137 256 141 259
rect 137 255 142 256
rect 105 249 111 254
rect 116 251 128 255
rect 132 251 133 255
rect 137 251 138 255
rect 105 247 107 249
rect 98 245 107 247
rect 137 250 142 251
rect 137 246 141 250
rect 98 241 111 245
rect 117 242 141 246
rect 91 240 95 241
rect 117 240 121 242
rect 33 235 37 236
rect 42 234 43 238
rect 47 234 66 238
rect 20 228 26 233
rect 104 233 105 237
rect 109 233 110 237
rect 146 238 150 267
rect 160 264 164 271
rect 160 263 165 264
rect 160 259 161 263
rect 168 263 172 284
rect 175 278 188 279
rect 175 274 178 278
rect 182 274 184 278
rect 175 273 188 274
rect 175 266 181 273
rect 191 267 195 284
rect 168 259 171 263
rect 175 259 176 263
rect 180 259 181 263
rect 185 259 186 263
rect 191 262 195 263
rect 160 258 165 259
rect 160 250 164 258
rect 180 254 186 259
rect 167 250 168 254
rect 172 250 186 254
rect 192 253 196 255
rect 117 235 121 236
rect 126 234 127 238
rect 131 234 150 238
rect 154 247 164 250
rect 154 235 157 247
rect 104 228 110 233
rect 160 241 164 247
rect 160 240 165 241
rect 160 236 161 240
rect 165 236 172 239
rect 160 233 172 236
rect 176 237 180 250
rect 192 246 196 249
rect 183 242 187 246
rect 191 242 196 246
rect 183 241 196 242
rect 176 233 190 237
rect 194 233 195 237
rect -73 224 -70 228
rect -66 224 -60 228
rect -56 224 8 228
rect 12 224 61 228
rect 65 224 92 228
rect 96 224 145 228
rect 149 224 162 228
rect 166 224 172 228
rect 176 227 200 228
rect 176 224 194 227
rect -87 221 194 224
rect -87 220 200 221
rect 17 218 61 220
rect 17 214 23 218
rect 27 214 51 218
rect 55 214 61 218
rect 21 206 27 214
rect 21 202 22 206
rect 26 202 27 206
rect 32 206 36 207
rect 41 206 47 214
rect 41 202 42 206
rect 46 202 47 206
rect 52 206 57 209
rect 56 202 57 206
rect 32 199 36 202
rect 52 201 57 202
rect 32 195 49 199
rect 21 183 25 193
rect 29 188 34 192
rect 45 191 49 195
rect 29 180 35 184
rect 39 180 42 184
rect -107 153 -102 173
rect 29 174 33 180
rect 45 176 49 187
rect 16 171 33 174
rect 37 172 49 176
rect 53 197 214 201
rect 37 168 41 172
rect 53 171 57 197
rect 223 175 227 284
rect 257 266 261 273
rect 257 265 262 266
rect 257 261 258 265
rect 265 265 269 286
rect 272 280 285 281
rect 272 276 275 280
rect 279 276 281 280
rect 272 275 285 276
rect 272 268 278 275
rect 288 269 292 286
rect 358 286 370 287
rect 374 287 454 290
rect 374 286 438 287
rect 335 275 347 281
rect 354 280 358 283
rect 442 286 454 287
rect 458 286 491 290
rect 495 286 505 290
rect 509 286 519 290
rect 523 289 586 290
rect 590 289 600 293
rect 604 289 614 293
rect 618 290 697 293
rect 618 289 681 290
rect 523 286 559 289
rect 368 277 390 281
rect 394 277 395 281
rect 410 280 431 281
rect 368 276 372 277
rect 354 275 358 276
rect 335 272 340 275
rect 335 271 336 272
rect 265 261 268 265
rect 272 261 273 265
rect 277 261 278 265
rect 282 261 283 265
rect 288 264 292 265
rect 327 268 336 271
rect 361 272 372 276
rect 410 276 424 280
rect 428 276 431 280
rect 410 275 431 276
rect 438 280 442 283
rect 452 277 474 281
rect 478 277 479 281
rect 452 276 456 277
rect 438 275 442 276
rect 361 268 365 272
rect 379 269 380 273
rect 384 269 395 273
rect 257 260 262 261
rect 257 252 261 260
rect 277 256 283 261
rect 264 252 265 256
rect 269 252 283 256
rect 289 254 293 257
rect 327 254 330 268
rect 335 267 340 268
rect 344 266 365 268
rect 257 243 261 248
rect 257 242 262 243
rect 257 238 258 242
rect 262 238 269 241
rect 257 235 269 238
rect 273 239 277 252
rect 336 262 344 263
rect 348 264 365 266
rect 336 259 348 262
rect 289 248 293 250
rect 280 244 284 248
rect 288 244 293 248
rect 280 243 293 244
rect 336 247 340 259
rect 361 257 365 264
rect 369 262 370 266
rect 374 265 375 266
rect 374 262 386 265
rect 369 261 386 262
rect 382 258 386 261
rect 382 257 387 258
rect 350 251 356 256
rect 361 253 373 257
rect 377 253 378 257
rect 382 253 383 257
rect 350 249 352 251
rect 343 247 352 249
rect 382 252 387 253
rect 391 253 395 269
rect 419 272 424 275
rect 419 268 420 272
rect 445 272 456 276
rect 445 268 449 272
rect 463 269 464 273
rect 468 269 481 273
rect 419 267 424 268
rect 428 266 449 268
rect 420 262 428 263
rect 432 264 449 266
rect 420 259 432 262
rect 382 248 386 252
rect 343 243 356 247
rect 362 244 386 248
rect 391 249 393 253
rect 336 242 340 243
rect 362 242 366 244
rect 273 235 287 239
rect 291 235 292 239
rect 349 235 350 239
rect 354 235 355 239
rect 391 240 395 249
rect 420 247 424 259
rect 445 257 449 264
rect 453 262 454 266
rect 458 265 459 266
rect 458 262 470 265
rect 453 261 470 262
rect 466 258 470 261
rect 466 257 471 258
rect 434 251 440 256
rect 445 253 457 257
rect 461 253 462 257
rect 466 253 467 257
rect 434 249 436 251
rect 427 247 436 249
rect 466 252 471 253
rect 466 248 470 252
rect 427 243 440 247
rect 446 244 470 248
rect 420 242 424 243
rect 446 242 450 244
rect 362 237 366 238
rect 371 236 372 240
rect 376 236 395 240
rect 349 230 355 235
rect 433 235 434 239
rect 438 235 439 239
rect 475 240 479 269
rect 489 266 493 273
rect 489 265 494 266
rect 489 261 490 265
rect 497 265 501 286
rect 504 280 517 281
rect 504 276 507 280
rect 511 276 513 280
rect 504 275 517 276
rect 504 268 510 275
rect 520 269 524 286
rect 497 261 500 265
rect 504 261 505 265
rect 509 261 510 265
rect 514 261 515 265
rect 520 264 524 265
rect 489 260 494 261
rect 489 252 493 260
rect 509 256 515 261
rect 496 252 497 256
rect 501 252 515 256
rect 521 255 525 257
rect 446 237 450 238
rect 455 236 456 240
rect 460 236 479 240
rect 483 249 493 252
rect 483 237 486 249
rect 433 230 439 235
rect 489 243 493 249
rect 489 242 494 243
rect 489 238 490 242
rect 494 238 501 241
rect 489 235 501 238
rect 505 239 509 252
rect 521 248 525 251
rect 512 244 516 248
rect 520 244 525 248
rect 512 243 525 244
rect 505 235 519 239
rect 523 235 524 239
rect 256 226 259 230
rect 263 226 269 230
rect 273 226 337 230
rect 341 226 390 230
rect 394 226 421 230
rect 425 226 474 230
rect 478 226 491 230
rect 495 226 501 230
rect 505 229 529 230
rect 505 226 521 229
rect 256 225 521 226
rect 241 223 521 225
rect 527 223 529 229
rect 241 222 529 223
rect 241 221 257 222
rect 346 220 390 222
rect 346 216 352 220
rect 356 216 380 220
rect 384 216 390 220
rect 350 208 356 216
rect 350 204 351 208
rect 355 204 356 208
rect 361 208 365 209
rect 370 208 376 216
rect 370 204 371 208
rect 375 204 376 208
rect 381 208 386 211
rect 385 204 386 208
rect 361 201 365 204
rect 381 203 386 204
rect 243 197 311 201
rect 361 197 378 201
rect 350 185 354 195
rect 358 190 363 194
rect 374 193 378 197
rect 358 182 364 186
rect 368 182 371 186
rect 52 170 57 171
rect 21 164 22 168
rect 26 164 41 168
rect 44 166 52 168
rect 56 166 57 170
rect 44 164 57 166
rect 39 158 40 161
rect 17 157 40 158
rect 44 158 45 161
rect 44 157 51 158
rect 17 154 51 157
rect 55 154 61 158
rect 17 153 61 154
rect 222 155 227 175
rect 358 176 362 182
rect 374 178 378 189
rect 345 173 362 176
rect 366 174 378 178
rect 382 197 386 203
rect 382 194 533 197
rect 537 194 538 197
rect 366 170 370 174
rect 382 173 386 194
rect 550 178 554 286
rect 584 269 588 276
rect 584 268 589 269
rect 584 264 585 268
rect 592 268 596 289
rect 599 283 612 284
rect 599 279 602 283
rect 606 279 608 283
rect 599 278 612 279
rect 599 271 605 278
rect 615 272 619 289
rect 685 289 697 290
rect 701 290 781 293
rect 701 289 765 290
rect 662 278 674 284
rect 681 283 685 286
rect 769 289 781 290
rect 785 289 818 293
rect 822 289 832 293
rect 836 289 846 293
rect 850 289 856 293
rect 695 280 717 284
rect 721 280 722 284
rect 735 283 758 284
rect 695 279 699 280
rect 735 279 751 283
rect 755 279 758 283
rect 681 278 685 279
rect 662 275 667 278
rect 662 274 663 275
rect 592 264 595 268
rect 599 264 600 268
rect 604 264 605 268
rect 609 264 610 268
rect 615 267 619 268
rect 584 263 589 264
rect 584 255 588 263
rect 604 259 610 264
rect 591 255 592 259
rect 596 255 610 259
rect 616 257 620 260
rect 584 246 588 251
rect 584 245 589 246
rect 584 241 585 245
rect 589 241 596 244
rect 584 238 596 241
rect 600 242 604 255
rect 616 251 620 253
rect 607 247 611 251
rect 615 247 620 251
rect 607 246 620 247
rect 600 238 614 242
rect 618 238 619 242
rect 643 240 647 269
rect 654 271 663 274
rect 688 275 699 279
rect 688 271 692 275
rect 706 272 707 276
rect 711 272 722 276
rect 654 257 657 271
rect 662 270 667 271
rect 671 269 692 271
rect 663 265 671 266
rect 675 267 692 269
rect 663 262 675 265
rect 663 250 667 262
rect 688 260 692 267
rect 696 265 697 269
rect 701 268 702 269
rect 701 265 713 268
rect 696 264 713 265
rect 709 261 713 264
rect 709 260 714 261
rect 677 254 683 259
rect 688 256 700 260
rect 704 256 705 260
rect 709 256 710 260
rect 677 252 679 254
rect 670 250 679 252
rect 709 255 714 256
rect 718 256 722 272
rect 709 251 713 255
rect 670 246 683 250
rect 689 247 713 251
rect 718 252 720 256
rect 663 245 667 246
rect 689 245 693 247
rect 643 236 644 240
rect 676 238 677 242
rect 681 238 682 242
rect 718 243 722 252
rect 689 240 693 241
rect 698 239 699 243
rect 703 239 722 243
rect 729 240 732 271
rect 676 233 682 238
rect 736 233 740 279
rect 746 278 758 279
rect 765 283 769 286
rect 779 280 801 284
rect 805 280 806 284
rect 779 279 783 280
rect 765 278 769 279
rect 746 275 751 278
rect 746 271 747 275
rect 772 275 783 279
rect 772 271 776 275
rect 790 272 791 276
rect 795 272 806 276
rect 746 270 751 271
rect 755 269 776 271
rect 747 265 755 266
rect 759 267 776 269
rect 747 262 759 265
rect 747 250 751 262
rect 772 260 776 267
rect 780 265 781 269
rect 785 268 786 269
rect 785 265 797 268
rect 780 264 797 265
rect 793 261 797 264
rect 793 260 798 261
rect 761 254 767 259
rect 772 256 784 260
rect 788 256 789 260
rect 793 256 794 260
rect 761 252 763 254
rect 754 250 763 252
rect 793 255 798 256
rect 793 251 797 255
rect 754 246 767 250
rect 773 247 797 251
rect 747 245 751 246
rect 773 245 777 247
rect 760 238 761 242
rect 765 238 766 242
rect 802 243 806 272
rect 816 269 820 276
rect 816 268 821 269
rect 816 264 817 268
rect 824 268 828 289
rect 831 283 844 284
rect 831 279 834 283
rect 838 279 840 283
rect 831 278 844 279
rect 831 271 837 278
rect 847 272 851 289
rect 824 264 827 268
rect 831 264 832 268
rect 836 264 837 268
rect 841 264 842 268
rect 847 267 851 268
rect 816 263 821 264
rect 816 255 820 263
rect 836 259 842 264
rect 823 255 824 259
rect 828 255 842 259
rect 848 258 852 260
rect 773 240 777 241
rect 782 239 783 243
rect 787 239 806 243
rect 810 252 820 255
rect 810 240 813 252
rect 760 233 766 238
rect 816 246 820 252
rect 816 245 821 246
rect 816 241 817 245
rect 821 241 828 244
rect 816 238 828 241
rect 832 242 836 255
rect 848 251 852 254
rect 839 247 843 251
rect 847 247 852 251
rect 839 246 852 247
rect 832 238 846 242
rect 850 238 851 242
rect 583 232 586 233
rect 581 229 586 232
rect 590 229 596 233
rect 600 229 664 233
rect 668 229 717 233
rect 721 229 748 233
rect 752 229 801 233
rect 805 229 818 233
rect 822 229 828 233
rect 832 229 856 233
rect 581 227 856 229
rect 568 225 856 227
rect 568 224 585 225
rect 568 223 584 224
rect 673 223 717 225
rect 673 219 679 223
rect 683 219 707 223
rect 711 219 717 223
rect 677 211 683 219
rect 677 207 678 211
rect 682 207 683 211
rect 688 211 692 212
rect 697 211 703 219
rect 697 207 698 211
rect 702 207 703 211
rect 708 211 713 214
rect 712 207 713 211
rect 569 194 636 197
rect 640 194 641 197
rect 381 172 386 173
rect 350 166 351 170
rect 355 166 370 170
rect 373 168 381 170
rect 385 168 386 172
rect 373 166 386 168
rect 368 160 369 163
rect 346 159 369 160
rect 373 160 374 163
rect 373 159 380 160
rect 346 156 380 159
rect 384 156 390 160
rect 346 155 390 156
rect -107 150 61 153
rect -107 149 21 150
rect 199 149 214 153
rect 18 146 21 149
rect 222 152 390 155
rect 549 158 554 178
rect 646 166 650 206
rect 688 204 692 207
rect 708 206 713 207
rect 688 200 705 204
rect 658 172 661 199
rect 677 188 681 198
rect 685 193 690 197
rect 701 196 705 200
rect 685 185 691 189
rect 695 185 698 189
rect 685 179 689 185
rect 701 181 705 192
rect 672 176 689 179
rect 693 177 705 181
rect 709 202 713 206
rect 709 199 721 202
rect 693 173 697 177
rect 709 176 713 199
rect 729 178 732 193
rect 708 175 713 176
rect 677 169 678 173
rect 682 169 697 173
rect 700 171 708 173
rect 712 171 713 175
rect 700 169 713 171
rect 695 163 696 166
rect 646 161 650 162
rect 673 162 696 163
rect 700 163 701 166
rect 728 165 733 178
rect 700 162 707 163
rect 673 159 707 162
rect 711 159 717 163
rect 673 158 717 159
rect 549 155 717 158
rect 549 154 673 155
rect 222 151 348 152
rect 678 151 681 155
rect 345 148 348 151
rect -107 142 199 146
rect -107 138 -71 142
rect -67 138 -57 142
rect -53 138 -43 142
rect -39 139 40 142
rect -39 138 24 139
rect -107 27 -103 138
rect -73 118 -69 125
rect -73 117 -68 118
rect -73 113 -72 117
rect -65 117 -61 138
rect -58 132 -45 133
rect -58 128 -55 132
rect -51 128 -49 132
rect -58 127 -45 128
rect -58 120 -52 127
rect -42 121 -38 138
rect 28 138 40 139
rect 44 139 124 142
rect 44 138 108 139
rect 5 127 17 133
rect 24 132 28 135
rect 112 138 124 139
rect 128 138 161 142
rect 165 138 175 142
rect 179 138 189 142
rect 193 138 199 142
rect 222 144 528 148
rect 222 140 258 144
rect 262 140 272 144
rect 276 140 286 144
rect 290 141 369 144
rect 290 140 353 141
rect 38 129 60 133
rect 64 129 65 133
rect 89 132 101 133
rect 77 129 94 132
rect 38 128 42 129
rect 24 127 28 128
rect 5 124 10 127
rect 5 123 6 124
rect -65 113 -62 117
rect -58 113 -57 117
rect -53 113 -52 117
rect -48 113 -47 117
rect -42 116 -38 117
rect -3 120 6 123
rect 31 124 42 128
rect 31 120 35 124
rect 49 121 50 125
rect 54 121 65 125
rect -73 112 -68 113
rect -73 104 -69 112
rect -53 108 -47 113
rect -66 104 -65 108
rect -61 104 -47 108
rect -41 106 -37 109
rect -3 106 0 120
rect 5 119 10 120
rect 14 118 35 120
rect -73 95 -69 100
rect -73 94 -68 95
rect -73 90 -72 94
rect -68 90 -61 93
rect -73 87 -61 90
rect -57 91 -53 104
rect 6 114 14 115
rect 18 116 35 118
rect 6 111 18 114
rect -41 100 -37 102
rect -50 96 -46 100
rect -42 96 -37 100
rect -50 95 -37 96
rect 6 99 10 111
rect 31 109 35 116
rect 39 114 40 118
rect 44 117 45 118
rect 44 114 56 117
rect 39 113 56 114
rect 52 110 56 113
rect 52 109 57 110
rect 20 103 26 108
rect 31 105 43 109
rect 47 105 48 109
rect 52 105 53 109
rect 20 101 22 103
rect 13 99 22 101
rect 52 104 57 105
rect 61 105 65 121
rect 52 100 56 104
rect 13 95 26 99
rect 32 96 56 100
rect 61 101 63 105
rect 6 94 10 95
rect 32 94 36 96
rect -57 87 -43 91
rect -39 87 -38 91
rect 19 87 20 91
rect 24 87 25 91
rect 61 92 65 101
rect 32 89 36 90
rect 41 88 42 92
rect 46 88 65 92
rect 77 89 80 129
rect 89 128 94 129
rect 98 128 101 132
rect 89 127 101 128
rect 108 132 112 135
rect 122 129 144 133
rect 148 129 149 133
rect 122 128 126 129
rect 108 127 112 128
rect 89 124 94 127
rect 89 120 90 124
rect 115 124 126 128
rect 115 120 119 124
rect 133 121 134 125
rect 138 121 149 125
rect 89 119 94 120
rect 98 118 119 120
rect 90 114 98 115
rect 102 116 119 118
rect 90 111 102 114
rect 90 99 94 111
rect 115 109 119 116
rect 123 114 124 118
rect 128 117 129 118
rect 128 114 140 117
rect 123 113 140 114
rect 136 110 140 113
rect 136 109 141 110
rect 104 103 110 108
rect 115 105 127 109
rect 131 105 132 109
rect 136 105 137 109
rect 104 101 106 103
rect 97 99 106 101
rect 136 104 141 105
rect 136 100 140 104
rect 97 95 110 99
rect 116 96 140 100
rect 90 94 94 95
rect 116 94 120 96
rect 19 82 25 87
rect 103 87 104 91
rect 108 87 109 91
rect 145 92 149 121
rect 159 118 163 125
rect 159 117 164 118
rect 159 113 160 117
rect 167 117 171 138
rect 174 132 187 133
rect 174 128 177 132
rect 181 128 183 132
rect 174 127 187 128
rect 174 120 180 127
rect 190 121 194 138
rect 167 113 170 117
rect 174 113 175 117
rect 179 113 180 117
rect 184 113 185 117
rect 190 116 194 117
rect 159 112 164 113
rect 159 104 163 112
rect 179 108 185 113
rect 166 104 167 108
rect 171 104 185 108
rect 191 107 195 109
rect 116 89 120 90
rect 125 88 126 92
rect 130 88 149 92
rect 153 101 163 104
rect 153 89 156 101
rect 103 82 109 87
rect 159 95 163 101
rect 159 94 164 95
rect 159 90 160 94
rect 164 90 171 93
rect 159 87 171 90
rect 175 91 179 104
rect 191 100 195 103
rect 182 96 186 100
rect 190 96 195 100
rect 182 95 195 96
rect 175 87 189 91
rect 193 87 194 91
rect -74 78 -71 82
rect -67 78 -61 82
rect -57 78 7 82
rect 11 78 60 82
rect 64 78 91 82
rect 95 78 144 82
rect 148 78 161 82
rect 165 78 171 82
rect 175 78 194 82
rect -74 75 194 78
rect -74 74 199 75
rect 16 72 60 74
rect 16 68 22 72
rect 26 68 50 72
rect 54 68 60 72
rect 20 60 26 68
rect 20 56 21 60
rect 25 56 26 60
rect 31 60 35 61
rect 40 60 46 68
rect 147 65 188 68
rect 40 56 41 60
rect 45 56 46 60
rect 51 60 56 63
rect 55 56 56 60
rect 31 53 35 56
rect 51 55 56 56
rect 31 49 48 53
rect 20 37 24 47
rect 28 42 33 46
rect 44 45 48 49
rect 28 34 34 38
rect 38 34 41 38
rect -108 7 -103 27
rect 28 28 32 34
rect 44 30 48 41
rect 15 25 32 28
rect 36 26 48 30
rect 36 22 40 26
rect 52 25 56 55
rect 144 47 167 50
rect 172 47 173 50
rect 51 24 56 25
rect 20 18 21 22
rect 25 18 40 22
rect 43 20 51 22
rect 55 20 56 24
rect 43 18 56 20
rect 38 12 39 15
rect 16 11 39 12
rect 43 12 44 15
rect 43 11 50 12
rect 16 8 50 11
rect 54 8 60 12
rect 16 7 60 8
rect -108 4 60 7
rect -108 3 16 4
rect 185 -36 188 65
rect 197 46 213 50
rect 222 29 226 140
rect 256 120 260 127
rect 256 119 261 120
rect 256 115 257 119
rect 264 119 268 140
rect 271 134 284 135
rect 271 130 274 134
rect 278 130 280 134
rect 271 129 284 130
rect 271 122 277 129
rect 287 123 291 140
rect 357 140 369 141
rect 373 141 453 144
rect 373 140 437 141
rect 334 129 346 135
rect 353 134 357 137
rect 441 140 453 141
rect 457 140 490 144
rect 494 140 504 144
rect 508 140 518 144
rect 522 140 528 144
rect 549 147 855 151
rect 549 143 585 147
rect 589 143 599 147
rect 603 143 613 147
rect 617 144 696 147
rect 617 143 680 144
rect 367 131 389 135
rect 393 131 394 135
rect 418 134 430 135
rect 367 130 371 131
rect 353 129 357 130
rect 334 126 339 129
rect 334 125 335 126
rect 264 115 267 119
rect 271 115 272 119
rect 276 115 277 119
rect 281 115 282 119
rect 287 118 291 119
rect 326 122 335 125
rect 360 126 371 130
rect 418 130 423 134
rect 427 130 430 134
rect 418 129 430 130
rect 437 134 441 137
rect 451 131 473 135
rect 477 131 478 135
rect 451 130 455 131
rect 437 129 441 130
rect 360 122 364 126
rect 378 123 379 127
rect 383 123 394 127
rect 256 114 261 115
rect 256 106 260 114
rect 276 110 282 115
rect 263 106 264 110
rect 268 106 282 110
rect 288 108 292 111
rect 256 97 260 102
rect 256 96 261 97
rect 256 92 257 96
rect 261 92 268 95
rect 256 89 268 92
rect 272 93 276 106
rect 288 102 292 104
rect 279 98 283 102
rect 287 98 292 102
rect 279 97 292 98
rect 272 89 286 93
rect 290 89 291 93
rect 316 91 319 111
rect 326 108 329 122
rect 334 121 339 122
rect 343 120 364 122
rect 335 116 343 117
rect 347 118 364 120
rect 335 113 347 116
rect 335 101 339 113
rect 360 111 364 118
rect 368 116 369 120
rect 373 119 374 120
rect 373 116 385 119
rect 368 115 385 116
rect 381 112 385 115
rect 381 111 386 112
rect 349 105 355 110
rect 360 107 372 111
rect 376 107 377 111
rect 381 107 382 111
rect 349 103 351 105
rect 342 101 351 103
rect 381 106 386 107
rect 390 107 394 123
rect 418 126 423 129
rect 418 122 419 126
rect 444 126 455 130
rect 444 122 448 126
rect 462 123 463 127
rect 467 123 478 127
rect 418 121 423 122
rect 427 120 448 122
rect 419 116 427 117
rect 431 118 448 120
rect 419 113 431 116
rect 381 102 385 106
rect 342 97 355 101
rect 361 98 385 102
rect 390 103 392 107
rect 335 96 339 97
rect 361 96 365 98
rect 348 89 349 93
rect 353 89 354 93
rect 390 94 394 103
rect 419 101 423 113
rect 444 111 448 118
rect 452 116 453 120
rect 457 119 458 120
rect 457 116 469 119
rect 452 115 469 116
rect 465 112 469 115
rect 465 111 470 112
rect 433 105 439 110
rect 444 107 456 111
rect 460 107 461 111
rect 465 107 466 111
rect 433 103 435 105
rect 426 101 435 103
rect 465 106 470 107
rect 465 102 469 106
rect 426 97 439 101
rect 445 98 469 102
rect 419 96 423 97
rect 445 96 449 98
rect 361 91 365 92
rect 370 90 371 94
rect 375 90 394 94
rect 348 84 354 89
rect 432 89 433 93
rect 437 89 438 93
rect 474 94 478 123
rect 488 120 492 127
rect 488 119 493 120
rect 488 115 489 119
rect 496 119 500 140
rect 503 134 516 135
rect 503 130 506 134
rect 510 130 512 134
rect 503 129 516 130
rect 503 122 509 129
rect 519 123 523 140
rect 496 115 499 119
rect 503 115 504 119
rect 508 115 509 119
rect 513 115 514 119
rect 519 118 523 119
rect 488 114 493 115
rect 488 106 492 114
rect 508 110 514 115
rect 495 106 496 110
rect 500 106 514 110
rect 520 109 524 111
rect 445 91 449 92
rect 454 90 455 94
rect 459 90 478 94
rect 482 103 492 106
rect 482 91 485 103
rect 432 84 438 89
rect 488 97 492 103
rect 488 96 493 97
rect 488 92 489 96
rect 493 92 500 95
rect 488 89 500 92
rect 504 93 508 106
rect 520 102 524 105
rect 511 98 515 102
rect 519 98 524 102
rect 511 97 524 98
rect 504 89 518 93
rect 522 89 523 93
rect 255 80 258 84
rect 262 80 268 84
rect 272 80 336 84
rect 340 80 389 84
rect 393 80 420 84
rect 424 80 473 84
rect 477 80 490 84
rect 494 80 500 84
rect 504 80 528 84
rect 236 77 521 80
rect 255 76 521 77
rect 525 76 528 80
rect 345 74 389 76
rect 345 70 351 74
rect 355 70 379 74
rect 383 70 389 74
rect 316 65 319 67
rect 349 62 355 70
rect 316 47 319 61
rect 349 58 350 62
rect 354 58 355 62
rect 360 62 364 63
rect 369 62 375 70
rect 369 58 370 62
rect 374 58 375 62
rect 380 62 385 65
rect 384 58 385 62
rect 360 55 364 58
rect 380 57 385 58
rect 360 51 377 55
rect 221 9 226 29
rect 288 43 316 46
rect 288 17 292 43
rect 349 39 353 49
rect 357 44 362 48
rect 373 47 377 51
rect 357 36 363 40
rect 367 36 370 40
rect 357 30 361 36
rect 373 32 377 43
rect 344 27 361 30
rect 365 28 377 32
rect 365 24 369 28
rect 381 27 385 57
rect 412 53 494 58
rect 549 32 553 143
rect 583 123 587 130
rect 583 122 588 123
rect 583 118 584 122
rect 591 122 595 143
rect 598 137 611 138
rect 598 133 601 137
rect 605 133 607 137
rect 598 132 611 133
rect 598 125 604 132
rect 614 126 618 143
rect 684 143 696 144
rect 700 144 780 147
rect 700 143 764 144
rect 661 132 673 138
rect 680 137 684 140
rect 768 143 780 144
rect 784 143 817 147
rect 821 143 831 147
rect 835 143 845 147
rect 849 143 855 147
rect 694 134 716 138
rect 720 134 721 138
rect 745 137 757 138
rect 694 133 698 134
rect 680 132 684 133
rect 661 129 666 132
rect 661 128 662 129
rect 591 118 594 122
rect 598 118 599 122
rect 603 118 604 122
rect 608 118 609 122
rect 614 121 618 122
rect 653 125 662 128
rect 687 129 698 133
rect 745 133 750 137
rect 754 133 757 137
rect 745 132 757 133
rect 764 137 768 140
rect 778 134 800 138
rect 804 134 805 138
rect 778 133 782 134
rect 764 132 768 133
rect 687 125 691 129
rect 705 126 706 130
rect 710 126 721 130
rect 583 117 588 118
rect 583 109 587 117
rect 603 113 609 118
rect 590 109 591 113
rect 595 109 609 113
rect 615 111 619 114
rect 653 111 656 125
rect 661 124 666 125
rect 670 123 691 125
rect 583 100 587 105
rect 583 99 588 100
rect 583 95 584 99
rect 588 95 595 98
rect 583 92 595 95
rect 599 96 603 109
rect 662 119 670 120
rect 674 121 691 123
rect 662 116 674 119
rect 615 105 619 107
rect 606 101 610 105
rect 614 101 619 105
rect 606 100 619 101
rect 662 104 666 116
rect 687 114 691 121
rect 695 119 696 123
rect 700 122 701 123
rect 700 119 712 122
rect 695 118 712 119
rect 708 115 712 118
rect 708 114 713 115
rect 676 108 682 113
rect 687 110 699 114
rect 703 110 704 114
rect 708 110 709 114
rect 676 106 678 108
rect 662 99 666 100
rect 669 104 678 106
rect 708 109 713 110
rect 717 110 721 126
rect 745 129 750 132
rect 745 125 746 129
rect 771 129 782 133
rect 771 125 775 129
rect 789 126 790 130
rect 794 126 805 130
rect 745 124 750 125
rect 754 123 775 125
rect 746 119 754 120
rect 758 121 775 123
rect 746 116 758 119
rect 708 105 712 109
rect 669 100 682 104
rect 688 101 712 105
rect 717 106 719 110
rect 599 92 613 96
rect 617 92 618 96
rect 669 95 672 100
rect 688 99 692 101
rect 658 91 672 95
rect 675 92 676 96
rect 680 92 681 96
rect 717 97 721 106
rect 746 104 750 116
rect 771 114 775 121
rect 779 119 780 123
rect 784 122 785 123
rect 784 119 796 122
rect 779 118 796 119
rect 792 115 796 118
rect 792 114 797 115
rect 760 108 766 113
rect 771 110 783 114
rect 787 110 788 114
rect 792 110 793 114
rect 760 106 762 108
rect 753 104 762 106
rect 792 109 797 110
rect 792 105 796 109
rect 753 100 766 104
rect 772 101 796 105
rect 746 99 750 100
rect 772 99 776 101
rect 688 94 692 95
rect 697 93 698 97
rect 702 93 721 97
rect 658 87 662 91
rect 675 87 681 92
rect 759 92 760 96
rect 764 92 765 96
rect 801 97 805 126
rect 815 123 819 130
rect 815 122 820 123
rect 815 118 816 122
rect 823 122 827 143
rect 830 137 843 138
rect 830 133 833 137
rect 837 133 839 137
rect 830 132 843 133
rect 830 125 836 132
rect 846 126 850 143
rect 823 118 826 122
rect 830 118 831 122
rect 835 118 836 122
rect 840 118 841 122
rect 846 121 850 122
rect 815 117 820 118
rect 815 109 819 117
rect 835 113 841 118
rect 822 109 823 113
rect 827 109 841 113
rect 847 112 851 114
rect 772 94 776 95
rect 781 93 782 97
rect 786 93 805 97
rect 809 106 819 109
rect 809 94 812 106
rect 759 87 765 92
rect 815 100 819 106
rect 815 99 820 100
rect 815 95 816 99
rect 820 95 827 98
rect 815 92 827 95
rect 831 96 835 109
rect 847 105 851 108
rect 838 101 842 105
rect 846 101 851 105
rect 838 100 851 101
rect 831 92 845 96
rect 849 92 850 96
rect 582 84 585 87
rect 581 83 585 84
rect 589 83 595 87
rect 599 83 663 87
rect 667 83 716 87
rect 720 83 747 87
rect 751 83 800 87
rect 804 83 817 87
rect 821 83 827 87
rect 831 83 855 87
rect 581 81 855 83
rect 562 80 855 81
rect 565 79 855 80
rect 565 78 584 79
rect 672 77 716 79
rect 672 73 678 77
rect 682 73 706 77
rect 710 73 716 77
rect 619 71 623 72
rect 563 53 592 58
rect 380 26 385 27
rect 349 20 350 24
rect 354 20 369 24
rect 372 22 380 24
rect 384 24 385 26
rect 384 22 389 24
rect 372 20 389 22
rect 367 14 368 17
rect 345 13 368 14
rect 372 14 373 17
rect 372 13 379 14
rect 345 10 379 13
rect 383 10 389 14
rect 345 9 389 10
rect 221 6 389 9
rect 548 12 553 32
rect 619 30 623 67
rect 676 65 682 73
rect 676 61 677 65
rect 681 61 682 65
rect 687 65 691 66
rect 696 65 702 73
rect 696 61 697 65
rect 701 61 702 65
rect 707 65 712 68
rect 711 61 712 65
rect 687 58 691 61
rect 707 60 712 61
rect 687 54 704 58
rect 676 42 680 52
rect 684 47 689 51
rect 700 50 704 54
rect 684 39 690 43
rect 694 39 697 43
rect 684 33 688 39
rect 700 35 704 46
rect 671 30 688 33
rect 692 31 704 35
rect 708 55 724 60
rect 692 27 696 31
rect 708 30 712 55
rect 707 29 712 30
rect 676 23 677 27
rect 681 23 696 27
rect 699 25 707 27
rect 711 25 712 29
rect 699 23 712 25
rect 694 17 695 20
rect 672 16 695 17
rect 699 17 700 20
rect 699 16 706 17
rect 672 13 706 16
rect 710 13 716 17
rect 672 12 716 13
rect 548 9 716 12
rect 548 8 672 9
rect 221 5 345 6
rect 334 -2 338 5
rect 217 -4 261 -2
rect 310 -4 354 -2
rect 397 -4 441 -2
rect 217 -6 441 -4
rect 217 -10 223 -6
rect 227 -7 316 -6
rect 227 -10 261 -7
rect 310 -10 316 -7
rect 320 -7 403 -6
rect 320 -10 354 -7
rect 397 -10 403 -7
rect 407 -10 441 -6
rect 231 -18 237 -10
rect 231 -22 232 -18
rect 236 -22 237 -18
rect 242 -16 246 -15
rect 251 -16 257 -10
rect 292 -16 303 -13
rect 251 -20 252 -16
rect 256 -20 257 -16
rect 221 -23 226 -22
rect 221 -27 222 -23
rect 242 -23 246 -20
rect 221 -30 226 -27
rect 221 -34 222 -30
rect 221 -35 226 -34
rect 229 -27 242 -25
rect 229 -29 246 -27
rect 253 -27 284 -23
rect 221 -36 225 -35
rect 185 -40 225 -36
rect 182 -52 212 -49
rect 221 -53 225 -40
rect 229 -40 233 -29
rect 244 -36 249 -32
rect 253 -36 257 -27
rect 236 -44 239 -40
rect 243 -44 250 -40
rect 229 -48 233 -44
rect 229 -52 241 -48
rect 245 -49 250 -44
rect 221 -54 226 -53
rect 221 -58 222 -54
rect 226 -58 233 -55
rect 221 -61 233 -58
rect 237 -56 241 -52
rect 244 -53 260 -49
rect 237 -60 252 -56
rect 256 -60 257 -56
rect 280 -60 284 -27
rect 300 -26 303 -16
rect 324 -18 330 -10
rect 324 -22 325 -18
rect 329 -22 330 -18
rect 335 -16 339 -15
rect 344 -16 350 -10
rect 344 -20 345 -16
rect 349 -20 350 -16
rect 411 -18 417 -10
rect 390 -19 406 -18
rect 314 -23 319 -22
rect 314 -26 315 -23
rect 300 -27 315 -26
rect 335 -23 339 -20
rect 300 -29 319 -27
rect 314 -30 319 -29
rect 314 -34 315 -30
rect 314 -35 319 -34
rect 322 -27 335 -25
rect 322 -29 339 -27
rect 314 -53 318 -35
rect 322 -40 326 -29
rect 346 -32 350 -23
rect 394 -23 406 -19
rect 411 -22 412 -18
rect 416 -22 417 -18
rect 422 -16 426 -15
rect 431 -16 437 -10
rect 431 -20 432 -16
rect 436 -20 437 -16
rect 394 -24 402 -23
rect 401 -27 402 -24
rect 422 -23 426 -20
rect 401 -30 406 -27
rect 337 -36 342 -32
rect 346 -36 357 -32
rect 401 -34 402 -30
rect 401 -35 406 -34
rect 409 -27 422 -25
rect 409 -29 426 -27
rect 329 -44 332 -40
rect 336 -44 343 -40
rect 322 -48 326 -44
rect 322 -52 334 -48
rect 314 -54 319 -53
rect 314 -58 315 -54
rect 319 -58 326 -55
rect 314 -61 326 -58
rect 330 -56 334 -52
rect 338 -49 343 -44
rect 338 -53 353 -49
rect 401 -53 405 -35
rect 409 -40 413 -29
rect 433 -32 437 -23
rect 424 -36 429 -32
rect 433 -36 446 -32
rect 416 -44 419 -40
rect 423 -44 430 -40
rect 409 -48 413 -44
rect 409 -52 421 -48
rect 401 -54 406 -53
rect 330 -60 345 -56
rect 349 -60 350 -56
rect 401 -58 402 -54
rect 406 -58 413 -55
rect 401 -61 413 -58
rect 417 -56 421 -52
rect 425 -50 430 -44
rect 425 -53 438 -50
rect 417 -60 432 -56
rect 436 -60 437 -56
rect 217 -70 223 -66
rect 227 -70 233 -66
rect 237 -70 261 -66
rect 310 -70 316 -66
rect 320 -70 326 -66
rect 330 -70 354 -66
rect 211 -71 354 -70
rect 397 -70 403 -66
rect 407 -70 413 -66
rect 417 -70 441 -66
rect 397 -71 441 -70
rect 211 -73 441 -71
rect 217 -74 261 -73
rect 310 -74 441 -73
<< metal2 >>
rect 206 410 308 413
rect 204 403 295 406
rect 205 396 276 399
rect -99 389 251 392
rect -27 370 2 374
rect -91 366 -24 370
rect -91 224 -86 366
rect -17 359 236 363
rect -76 301 -72 352
rect -17 324 -12 359
rect 231 355 235 359
rect 1 346 2 349
rect 6 346 90 349
rect 94 346 183 349
rect 87 328 231 331
rect -18 320 -6 324
rect 87 324 90 328
rect -1 320 10 324
rect 139 319 140 322
rect -77 299 -72 301
rect -77 263 -73 299
rect 67 298 115 301
rect 67 297 124 298
rect 112 294 124 297
rect 137 288 140 319
rect 180 314 183 320
rect 180 311 231 314
rect 246 311 251 389
rect 273 324 276 396
rect 292 335 295 403
rect 304 393 308 410
rect 304 357 307 393
rect 366 345 370 379
rect 408 360 656 364
rect 408 356 412 360
rect 416 348 461 349
rect 465 348 554 351
rect 380 347 383 348
rect 378 344 383 347
rect 416 347 554 348
rect 558 347 641 351
rect 416 346 464 347
rect 416 344 419 346
rect 378 341 419 344
rect 378 311 383 341
rect 413 330 560 333
rect 557 326 560 330
rect 461 322 465 325
rect 461 314 464 322
rect 413 311 464 314
rect 557 322 558 326
rect 575 324 594 328
rect 652 326 656 360
rect 638 322 646 326
rect 651 324 656 326
rect 651 322 878 324
rect 246 306 383 311
rect 248 305 257 306
rect 458 303 461 311
rect 385 300 396 302
rect 458 300 472 303
rect 385 299 390 300
rect 166 296 390 299
rect 394 296 396 300
rect 166 295 396 296
rect 496 294 499 321
rect 558 312 561 322
rect 652 321 878 322
rect 665 320 878 321
rect 864 312 868 313
rect 558 308 868 312
rect 511 300 570 303
rect 401 291 499 294
rect 598 300 860 303
rect 584 296 588 299
rect 584 293 651 296
rect 89 287 142 288
rect 7 284 142 287
rect 401 286 405 291
rect 7 278 10 284
rect -44 275 21 278
rect -77 259 -36 263
rect -40 252 -36 259
rect -87 220 -86 224
rect -79 250 -76 251
rect -79 247 -72 250
rect -79 182 -76 247
rect -36 248 -3 251
rect 17 251 20 275
rect 99 275 184 278
rect 188 275 209 278
rect 285 277 350 280
rect 68 247 101 250
rect 81 243 84 247
rect 193 243 196 249
rect 81 240 196 243
rect 157 231 158 234
rect 155 183 158 231
rect 206 225 209 275
rect 346 274 350 277
rect 401 274 404 286
rect 647 283 651 293
rect 408 280 428 282
rect 408 279 424 280
rect 408 275 409 279
rect 413 276 424 279
rect 428 277 513 280
rect 612 280 677 283
rect 413 275 428 276
rect 408 274 416 275
rect 346 271 404 274
rect 250 249 257 252
rect 200 221 234 225
rect 194 220 234 221
rect -79 179 15 182
rect 25 180 168 183
rect 12 175 15 179
rect 163 149 194 153
rect 144 148 168 149
rect 101 145 168 148
rect 101 144 104 145
rect 45 141 104 144
rect 45 132 49 141
rect -45 129 49 132
rect -80 101 -73 104
rect -80 36 -77 101
rect -37 102 -4 105
rect 16 105 19 129
rect 98 129 183 132
rect -23 67 -20 102
rect 67 101 100 104
rect 80 97 83 101
rect 192 97 195 103
rect 80 94 195 97
rect 156 85 157 88
rect 77 69 80 85
rect -23 63 70 67
rect 76 66 143 69
rect 65 50 70 63
rect 65 46 138 50
rect 154 37 157 85
rect 207 81 210 220
rect 218 197 239 201
rect 250 184 253 249
rect 293 250 326 253
rect 346 253 349 271
rect 485 269 643 272
rect 311 201 315 250
rect 397 249 430 252
rect 410 245 413 249
rect 522 245 525 251
rect 410 242 525 245
rect 577 252 584 255
rect 486 233 487 236
rect 484 185 487 233
rect 527 223 561 227
rect 521 222 561 223
rect 537 194 565 197
rect 577 187 580 252
rect 620 253 653 256
rect 673 256 676 280
rect 755 280 840 283
rect 732 272 806 274
rect 732 271 810 272
rect 636 198 640 253
rect 724 252 757 255
rect 737 248 740 252
rect 849 248 852 254
rect 737 245 852 248
rect 645 211 648 236
rect 813 236 814 239
rect 662 199 721 202
rect 729 198 733 236
rect 811 188 814 236
rect 250 181 344 184
rect 354 182 497 185
rect 577 184 671 187
rect 681 185 824 188
rect 341 177 344 181
rect 668 180 671 184
rect 639 173 659 176
rect 639 171 642 173
rect 399 168 642 171
rect 656 172 659 173
rect 719 173 767 176
rect 656 168 658 172
rect 662 168 663 171
rect 399 152 402 168
rect 719 164 722 173
rect 650 162 722 164
rect 646 161 722 162
rect 728 155 733 158
rect 219 149 402 152
rect 428 151 733 155
rect 428 150 551 151
rect 429 134 434 150
rect 761 137 764 173
rect 284 131 349 134
rect 316 115 319 131
rect 249 103 256 106
rect 202 80 232 81
rect 202 75 231 80
rect 172 46 192 50
rect -80 33 14 36
rect 24 34 167 37
rect 11 29 14 33
rect 203 -40 209 75
rect 230 50 234 51
rect 218 46 234 50
rect 230 25 234 46
rect 249 38 252 103
rect 292 104 325 107
rect 345 107 348 131
rect 427 131 512 134
rect 611 134 676 137
rect 307 57 310 104
rect 396 103 429 106
rect 409 99 412 103
rect 521 99 524 105
rect 409 96 524 99
rect 576 106 583 109
rect 316 91 319 92
rect 485 87 486 90
rect 316 65 319 87
rect 307 53 406 57
rect 483 39 486 87
rect 525 77 561 80
rect 499 53 558 58
rect 576 41 579 106
rect 619 107 652 110
rect 672 110 675 134
rect 754 134 839 137
rect 639 71 643 107
rect 723 106 756 109
rect 736 102 739 106
rect 848 102 851 108
rect 736 99 851 102
rect 812 90 813 93
rect 623 67 643 71
rect 639 66 643 67
rect 597 55 724 58
rect 730 55 731 58
rect 597 54 731 55
rect 810 42 813 90
rect 249 35 343 38
rect 353 36 496 39
rect 576 38 670 41
rect 680 39 823 42
rect 340 31 343 35
rect 667 34 670 38
rect 619 30 623 31
rect 230 21 307 25
rect 304 17 307 21
rect 387 20 389 25
rect 387 17 392 20
rect 288 -12 292 13
rect 304 13 392 17
rect 304 12 307 13
rect 619 -19 623 26
rect 857 20 860 300
rect 394 -22 623 -19
rect 394 -23 619 -22
rect 856 -32 860 20
rect 361 -36 395 -32
rect 450 -35 860 -32
rect 856 -36 860 -35
rect 391 -40 395 -36
rect 203 -68 206 -40
rect 391 -43 460 -40
rect 457 -47 460 -43
rect 864 -47 868 308
rect 217 -52 260 -49
rect 265 -53 353 -49
rect 358 -53 438 -50
rect 457 -51 868 -47
rect 875 -61 878 320
rect 284 -64 878 -61
rect 203 -75 204 -68
<< metal3 >>
rect 389 300 414 302
rect 389 296 390 300
rect 394 296 414 300
rect 389 295 395 296
rect 408 281 414 296
rect 408 279 415 281
rect 408 275 409 279
rect 413 275 415 279
rect 408 274 415 275
<< ntransistor >>
rect 13 347 15 358
rect 20 347 22 358
rect 33 347 35 356
rect 100 347 102 358
rect 107 347 109 358
rect 120 347 122 356
rect 193 347 195 358
rect 200 347 202 358
rect 213 347 215 356
rect 433 349 435 358
rect 446 349 448 360
rect 453 349 455 360
rect 526 349 528 358
rect 539 349 541 360
rect 546 349 548 360
rect 613 349 615 358
rect 626 349 628 360
rect 633 349 635 360
rect -65 235 -63 241
rect -53 229 -51 238
rect -46 229 -44 238
rect 13 237 15 246
rect 29 232 31 241
rect 39 232 41 241
rect 49 229 51 241
rect 56 229 58 241
rect 97 237 99 246
rect 113 232 115 241
rect 123 232 125 241
rect 133 229 135 241
rect 140 229 142 241
rect 167 235 169 241
rect 179 229 181 238
rect 186 229 188 238
rect 264 237 266 243
rect 276 231 278 240
rect 283 231 285 240
rect 342 239 344 248
rect 358 234 360 243
rect 368 234 370 243
rect 378 231 380 243
rect 385 231 387 243
rect 426 239 428 248
rect 442 234 444 243
rect 452 234 454 243
rect 462 231 464 243
rect 469 231 471 243
rect 496 237 498 243
rect 591 240 593 246
rect 508 231 510 240
rect 515 231 517 240
rect 603 234 605 243
rect 610 234 612 243
rect 669 242 671 251
rect 685 237 687 246
rect 695 237 697 246
rect 705 234 707 246
rect 712 234 714 246
rect 753 242 755 251
rect 769 237 771 246
rect 779 237 781 246
rect 789 234 791 246
rect 796 234 798 246
rect 823 240 825 246
rect 835 234 837 243
rect 842 234 844 243
rect 28 201 30 207
rect 38 201 40 207
rect 48 201 50 207
rect 357 203 359 209
rect 367 203 369 209
rect 377 203 379 209
rect 684 206 686 212
rect 694 206 696 212
rect 704 206 706 212
rect -66 89 -64 95
rect -54 83 -52 92
rect -47 83 -45 92
rect 12 91 14 100
rect 28 86 30 95
rect 38 86 40 95
rect 48 83 50 95
rect 55 83 57 95
rect 96 91 98 100
rect 112 86 114 95
rect 122 86 124 95
rect 132 83 134 95
rect 139 83 141 95
rect 166 89 168 95
rect 178 83 180 92
rect 185 83 187 92
rect 263 91 265 97
rect 275 85 277 94
rect 282 85 284 94
rect 341 93 343 102
rect 357 88 359 97
rect 367 88 369 97
rect 377 85 379 97
rect 384 85 386 97
rect 425 93 427 102
rect 441 88 443 97
rect 451 88 453 97
rect 461 85 463 97
rect 468 85 470 97
rect 495 91 497 97
rect 590 94 592 100
rect 507 85 509 94
rect 514 85 516 94
rect 602 88 604 97
rect 609 88 611 97
rect 668 96 670 105
rect 684 91 686 100
rect 694 91 696 100
rect 704 88 706 100
rect 711 88 713 100
rect 752 96 754 105
rect 768 91 770 100
rect 778 91 780 100
rect 788 88 790 100
rect 795 88 797 100
rect 822 94 824 100
rect 834 88 836 97
rect 841 88 843 97
rect 27 55 29 61
rect 37 55 39 61
rect 47 55 49 61
rect 356 57 358 63
rect 366 57 368 63
rect 376 57 378 63
rect 683 60 685 66
rect 693 60 695 66
rect 703 60 705 66
rect 228 -59 230 -50
rect 241 -61 243 -50
rect 248 -61 250 -50
rect 321 -59 323 -50
rect 334 -61 336 -50
rect 341 -61 343 -50
rect 408 -59 410 -50
rect 421 -61 423 -50
rect 428 -61 430 -50
<< ptransistor >>
rect 13 312 15 325
rect 23 312 25 325
rect 33 314 35 332
rect 100 312 102 325
rect 110 312 112 325
rect 120 314 122 332
rect 193 312 195 325
rect 203 312 205 325
rect 213 314 215 332
rect 433 316 435 334
rect 443 314 445 327
rect 453 314 455 327
rect 526 316 528 334
rect 536 314 538 327
rect 546 314 548 327
rect 613 316 615 334
rect 623 314 625 327
rect 633 314 635 327
rect -65 258 -63 270
rect -55 258 -53 268
rect -45 258 -43 268
rect 21 259 23 286
rect 37 259 39 277
rect 47 259 49 277
rect 57 259 59 286
rect 105 259 107 286
rect 121 259 123 277
rect 131 259 133 277
rect 141 259 143 286
rect 167 258 169 270
rect 177 258 179 268
rect 187 258 189 268
rect 264 260 266 272
rect 274 260 276 270
rect 284 260 286 270
rect 350 261 352 288
rect 366 261 368 279
rect 376 261 378 279
rect 386 261 388 288
rect 434 261 436 288
rect 450 261 452 279
rect 460 261 462 279
rect 470 261 472 288
rect 496 260 498 272
rect 506 260 508 270
rect 516 260 518 270
rect 591 263 593 275
rect 601 263 603 273
rect 611 263 613 273
rect 677 264 679 291
rect 693 264 695 282
rect 703 264 705 282
rect 713 264 715 291
rect 761 264 763 291
rect 777 264 779 282
rect 787 264 789 282
rect 797 264 799 291
rect 823 263 825 275
rect 833 263 835 273
rect 843 263 845 273
rect 28 156 30 174
rect 35 156 37 174
rect 48 165 50 177
rect 357 158 359 176
rect 364 158 366 176
rect 377 167 379 179
rect 684 161 686 179
rect 691 161 693 179
rect 704 170 706 182
rect -66 112 -64 124
rect -56 112 -54 122
rect -46 112 -44 122
rect 20 113 22 140
rect 36 113 38 131
rect 46 113 48 131
rect 56 113 58 140
rect 104 113 106 140
rect 120 113 122 131
rect 130 113 132 131
rect 140 113 142 140
rect 166 112 168 124
rect 176 112 178 122
rect 186 112 188 122
rect 263 114 265 126
rect 273 114 275 124
rect 283 114 285 124
rect 349 115 351 142
rect 365 115 367 133
rect 375 115 377 133
rect 385 115 387 142
rect 433 115 435 142
rect 449 115 451 133
rect 459 115 461 133
rect 469 115 471 142
rect 495 114 497 126
rect 505 114 507 124
rect 515 114 517 124
rect 590 117 592 129
rect 600 117 602 127
rect 610 117 612 127
rect 676 118 678 145
rect 692 118 694 136
rect 702 118 704 136
rect 712 118 714 145
rect 760 118 762 145
rect 776 118 778 136
rect 786 118 788 136
rect 796 118 798 145
rect 822 117 824 129
rect 832 117 834 127
rect 842 117 844 127
rect 27 10 29 28
rect 34 10 36 28
rect 47 19 49 31
rect 356 12 358 30
rect 363 12 365 30
rect 376 21 378 33
rect 683 15 685 33
rect 690 15 692 33
rect 703 24 705 36
rect 228 -35 230 -17
rect 238 -28 240 -15
rect 248 -28 250 -15
rect 321 -35 323 -17
rect 331 -28 333 -15
rect 341 -28 343 -15
rect 408 -35 410 -17
rect 418 -28 420 -15
rect 428 -28 430 -15
<< polycontact >>
rect 20 337 24 341
rect 30 337 34 341
rect 10 329 14 333
rect 107 337 111 341
rect 117 337 121 341
rect 97 329 101 333
rect 200 337 204 341
rect 210 337 214 341
rect 190 329 194 333
rect 434 339 438 343
rect 444 339 448 343
rect 527 339 531 343
rect 537 339 541 343
rect 454 331 458 335
rect 614 339 618 343
rect 624 339 628 343
rect 547 331 551 335
rect 634 331 638 335
rect -54 274 -50 278
rect 7 266 11 270
rect -64 250 -60 254
rect 91 266 95 270
rect 44 251 48 255
rect 54 251 58 255
rect 178 274 182 278
rect 275 276 279 280
rect 336 268 340 272
rect -45 242 -41 246
rect 23 245 27 249
rect 128 251 132 255
rect 138 251 142 255
rect 168 250 172 254
rect 107 245 111 249
rect 265 252 269 256
rect 187 242 191 246
rect 420 268 424 272
rect 373 253 377 257
rect 383 253 387 257
rect 507 276 511 280
rect 602 279 606 283
rect 663 271 667 275
rect 284 244 288 248
rect 352 247 356 251
rect 457 253 461 257
rect 467 253 471 257
rect 497 252 501 256
rect 436 247 440 251
rect 592 255 596 259
rect 516 244 520 248
rect 747 271 751 275
rect 700 256 704 260
rect 710 256 714 260
rect 834 279 838 283
rect 611 247 615 251
rect 679 250 683 254
rect 784 256 788 260
rect 794 256 798 260
rect 824 255 828 259
rect 763 250 767 254
rect 843 247 847 251
rect 25 188 29 192
rect 37 188 41 192
rect 45 187 49 191
rect 354 190 358 194
rect 366 190 370 194
rect 35 180 39 184
rect 374 189 378 193
rect 681 193 685 197
rect 693 193 697 197
rect 364 182 368 186
rect 701 192 705 196
rect 691 185 695 189
rect -55 128 -51 132
rect 6 120 10 124
rect -65 104 -61 108
rect 90 120 94 124
rect 43 105 47 109
rect 53 105 57 109
rect 177 128 181 132
rect 274 130 278 134
rect 335 122 339 126
rect -46 96 -42 100
rect 22 99 26 103
rect 127 105 131 109
rect 137 105 141 109
rect 167 104 171 108
rect 106 99 110 103
rect 264 106 268 110
rect 186 96 190 100
rect 419 122 423 126
rect 372 107 376 111
rect 382 107 386 111
rect 506 130 510 134
rect 601 133 605 137
rect 662 125 666 129
rect 283 98 287 102
rect 351 101 355 105
rect 456 107 460 111
rect 466 107 470 111
rect 496 106 500 110
rect 435 101 439 105
rect 591 109 595 113
rect 515 98 519 102
rect 746 125 750 129
rect 699 110 703 114
rect 709 110 713 114
rect 833 133 837 137
rect 610 101 614 105
rect 678 104 682 108
rect 783 110 787 114
rect 793 110 797 114
rect 823 109 827 113
rect 762 104 766 108
rect 842 101 846 105
rect 24 42 28 46
rect 36 42 40 46
rect 44 41 48 45
rect 353 44 357 48
rect 365 44 369 48
rect 34 34 38 38
rect 373 43 377 47
rect 680 47 684 51
rect 692 47 696 51
rect 363 36 367 40
rect 700 46 704 50
rect 690 39 694 43
rect 249 -36 253 -32
rect 229 -44 233 -40
rect 239 -44 243 -40
rect 342 -36 346 -32
rect 322 -44 326 -40
rect 332 -44 336 -40
rect 429 -36 433 -32
rect 409 -44 413 -40
rect 419 -44 423 -40
<< ndcontact >>
rect 26 363 30 367
rect 113 363 117 367
rect 7 353 11 357
rect 206 363 210 367
rect 37 351 41 355
rect 94 353 98 357
rect 438 365 442 369
rect 124 351 128 355
rect 187 353 191 357
rect 531 365 535 369
rect 217 351 221 355
rect 427 353 431 357
rect 457 355 461 359
rect 618 365 622 369
rect 520 353 524 357
rect 550 355 554 359
rect 607 353 611 357
rect 637 355 641 359
rect -71 236 -67 240
rect 7 241 11 245
rect 91 241 95 245
rect -42 233 -38 237
rect 21 233 25 237
rect 33 236 37 240
rect 43 234 47 238
rect -60 224 -56 228
rect 105 233 109 237
rect 117 236 121 240
rect 127 234 131 238
rect 61 224 65 228
rect 161 236 165 240
rect 258 238 262 242
rect 336 243 340 247
rect 190 233 194 237
rect 420 243 424 247
rect 287 235 291 239
rect 350 235 354 239
rect 362 238 366 242
rect 372 236 376 240
rect 145 224 149 228
rect 172 224 176 228
rect 269 226 273 230
rect 434 235 438 239
rect 446 238 450 242
rect 456 236 460 240
rect 390 226 394 230
rect 490 238 494 242
rect 585 241 589 245
rect 663 246 667 250
rect 519 235 523 239
rect 747 246 751 250
rect 614 238 618 242
rect 677 238 681 242
rect 689 241 693 245
rect 699 239 703 243
rect 474 226 478 230
rect 501 226 505 230
rect 596 229 600 233
rect 761 238 765 242
rect 773 241 777 245
rect 783 239 787 243
rect 717 229 721 233
rect 817 241 821 245
rect 846 238 850 242
rect 801 229 805 233
rect 828 229 832 233
rect 22 202 26 206
rect 32 202 36 206
rect 42 202 46 206
rect 52 202 56 206
rect 351 204 355 208
rect 361 204 365 208
rect 371 204 375 208
rect 381 204 385 208
rect 678 207 682 211
rect 688 207 692 211
rect 698 207 702 211
rect 708 207 712 211
rect -72 90 -68 94
rect 6 95 10 99
rect 90 95 94 99
rect -43 87 -39 91
rect 20 87 24 91
rect 32 90 36 94
rect 42 88 46 92
rect -61 78 -57 82
rect 104 87 108 91
rect 116 90 120 94
rect 126 88 130 92
rect 60 78 64 82
rect 160 90 164 94
rect 257 92 261 96
rect 335 97 339 101
rect 189 87 193 91
rect 419 97 423 101
rect 286 89 290 93
rect 349 89 353 93
rect 361 92 365 96
rect 371 90 375 94
rect 144 78 148 82
rect 171 78 175 82
rect 268 80 272 84
rect 433 89 437 93
rect 445 92 449 96
rect 455 90 459 94
rect 389 80 393 84
rect 489 92 493 96
rect 584 95 588 99
rect 662 100 666 104
rect 518 89 522 93
rect 746 100 750 104
rect 613 92 617 96
rect 676 92 680 96
rect 688 95 692 99
rect 698 93 702 97
rect 473 80 477 84
rect 500 80 504 84
rect 595 83 599 87
rect 760 92 764 96
rect 772 95 776 99
rect 782 93 786 97
rect 716 83 720 87
rect 816 95 820 99
rect 845 92 849 96
rect 800 83 804 87
rect 827 83 831 87
rect 21 56 25 60
rect 31 56 35 60
rect 41 56 45 60
rect 51 56 55 60
rect 350 58 354 62
rect 360 58 364 62
rect 370 58 374 62
rect 380 58 384 62
rect 677 61 681 65
rect 687 61 691 65
rect 697 61 701 65
rect 707 61 711 65
rect 222 -58 226 -54
rect 252 -60 256 -56
rect 315 -58 319 -54
rect 345 -60 349 -56
rect 402 -58 406 -54
rect 233 -70 237 -66
rect 432 -60 436 -56
rect 326 -70 330 -66
rect 413 -70 417 -66
<< pdcontact >>
rect 7 313 11 317
rect 17 320 21 324
rect 17 313 21 317
rect 27 315 31 319
rect 37 327 41 331
rect 37 320 41 324
rect 94 313 98 317
rect 104 320 108 324
rect 104 313 108 317
rect 114 315 118 319
rect 124 327 128 331
rect 124 320 128 324
rect 187 313 191 317
rect 197 320 201 324
rect 197 313 201 317
rect 207 315 211 319
rect 217 327 221 331
rect 217 320 221 324
rect 427 329 431 333
rect 427 322 431 326
rect 520 329 524 333
rect 437 317 441 321
rect 447 322 451 326
rect 447 315 451 319
rect 520 322 524 326
rect 457 315 461 319
rect 607 329 611 333
rect 530 317 534 321
rect 540 322 544 326
rect 540 315 544 319
rect 607 322 611 326
rect 550 315 554 319
rect 617 317 621 321
rect 627 322 631 326
rect 627 315 631 319
rect 637 315 641 319
rect -71 259 -67 263
rect -61 259 -57 263
rect -51 259 -47 263
rect -41 263 -37 267
rect 15 260 19 264
rect 25 281 29 285
rect 25 274 29 278
rect 41 260 45 264
rect 51 267 55 271
rect 61 275 65 279
rect 99 260 103 264
rect 109 281 113 285
rect 109 274 113 278
rect 125 260 129 264
rect 135 267 139 271
rect 145 275 149 279
rect 161 259 165 263
rect 171 259 175 263
rect 181 259 185 263
rect 191 263 195 267
rect 258 261 262 265
rect 268 261 272 265
rect 278 261 282 265
rect 288 265 292 269
rect 344 262 348 266
rect 354 283 358 287
rect 354 276 358 280
rect 370 262 374 266
rect 380 269 384 273
rect 390 277 394 281
rect 428 262 432 266
rect 438 283 442 287
rect 438 276 442 280
rect 454 262 458 266
rect 464 269 468 273
rect 474 277 478 281
rect 490 261 494 265
rect 500 261 504 265
rect 510 261 514 265
rect 520 265 524 269
rect 585 264 589 268
rect 595 264 599 268
rect 605 264 609 268
rect 615 268 619 272
rect 671 265 675 269
rect 681 286 685 290
rect 681 279 685 283
rect 697 265 701 269
rect 707 272 711 276
rect 717 280 721 284
rect 755 265 759 269
rect 765 286 769 290
rect 765 279 769 283
rect 781 265 785 269
rect 791 272 795 276
rect 801 280 805 284
rect 817 264 821 268
rect 827 264 831 268
rect 837 264 841 268
rect 847 268 851 272
rect 22 164 26 168
rect 52 166 56 170
rect 351 166 355 170
rect 40 157 44 161
rect 381 168 385 172
rect 678 169 682 173
rect 369 159 373 163
rect 708 171 712 175
rect 696 162 700 166
rect -72 113 -68 117
rect -62 113 -58 117
rect -52 113 -48 117
rect -42 117 -38 121
rect 14 114 18 118
rect 24 135 28 139
rect 24 128 28 132
rect 40 114 44 118
rect 50 121 54 125
rect 60 129 64 133
rect 98 114 102 118
rect 108 135 112 139
rect 108 128 112 132
rect 124 114 128 118
rect 134 121 138 125
rect 144 129 148 133
rect 160 113 164 117
rect 170 113 174 117
rect 180 113 184 117
rect 190 117 194 121
rect 257 115 261 119
rect 267 115 271 119
rect 277 115 281 119
rect 287 119 291 123
rect 343 116 347 120
rect 353 137 357 141
rect 353 130 357 134
rect 369 116 373 120
rect 379 123 383 127
rect 389 131 393 135
rect 427 116 431 120
rect 437 137 441 141
rect 437 130 441 134
rect 453 116 457 120
rect 463 123 467 127
rect 473 131 477 135
rect 489 115 493 119
rect 499 115 503 119
rect 509 115 513 119
rect 519 119 523 123
rect 584 118 588 122
rect 594 118 598 122
rect 604 118 608 122
rect 614 122 618 126
rect 670 119 674 123
rect 680 140 684 144
rect 680 133 684 137
rect 696 119 700 123
rect 706 126 710 130
rect 716 134 720 138
rect 754 119 758 123
rect 764 140 768 144
rect 764 133 768 137
rect 780 119 784 123
rect 790 126 794 130
rect 800 134 804 138
rect 816 118 820 122
rect 826 118 830 122
rect 836 118 840 122
rect 846 122 850 126
rect 21 18 25 22
rect 51 20 55 24
rect 350 20 354 24
rect 39 11 43 15
rect 380 22 384 26
rect 677 23 681 27
rect 368 13 372 17
rect 707 25 711 29
rect 695 16 699 20
rect 222 -27 226 -23
rect 222 -34 226 -30
rect 232 -22 236 -18
rect 242 -20 246 -16
rect 242 -27 246 -23
rect 252 -20 256 -16
rect 315 -27 319 -23
rect 315 -34 319 -30
rect 325 -22 329 -18
rect 335 -20 339 -16
rect 335 -27 339 -23
rect 345 -20 349 -16
rect 402 -27 406 -23
rect 402 -34 406 -30
rect 412 -22 416 -18
rect 422 -20 426 -16
rect 422 -27 426 -23
rect 432 -20 436 -16
<< m2contact >>
rect 366 379 371 385
rect 2 370 7 375
rect -76 352 -71 358
rect 2 346 6 350
rect -6 320 -1 325
rect 90 346 94 350
rect 86 320 90 324
rect 183 346 187 350
rect 231 351 235 355
rect 304 351 310 357
rect 407 351 412 356
rect 135 319 139 323
rect 179 320 183 324
rect 365 340 370 345
rect 231 328 235 332
rect 292 329 298 335
rect 461 348 465 352
rect 408 328 413 333
rect 273 318 279 324
rect 465 322 469 326
rect 231 311 235 315
rect 409 311 413 315
rect 496 321 500 326
rect 554 347 558 351
rect 641 347 645 351
rect 558 322 562 326
rect 571 324 575 328
rect 124 294 128 298
rect 161 295 166 299
rect 472 300 477 305
rect 507 300 511 305
rect 570 300 574 304
rect 584 299 588 303
rect 594 324 598 328
rect 646 322 651 326
rect 594 300 598 304
rect -48 274 -44 278
rect 95 274 99 278
rect -72 246 -68 250
rect -40 248 -36 252
rect -3 248 1 252
rect 17 247 21 251
rect 64 247 68 251
rect 101 247 105 251
rect 184 274 188 278
rect 153 231 157 235
rect 192 249 196 253
rect -91 220 -87 224
rect 194 221 200 227
rect 21 179 25 183
rect 12 171 16 175
rect 214 197 218 201
rect 281 276 285 280
rect 424 276 428 280
rect 257 248 261 252
rect 289 250 293 254
rect 326 250 330 254
rect 346 249 350 253
rect 481 269 485 273
rect 393 249 397 253
rect 430 249 434 253
rect 513 276 517 280
rect 482 233 486 237
rect 521 251 525 255
rect 234 220 241 227
rect 521 223 527 229
rect 239 197 243 201
rect 311 197 315 201
rect 350 181 354 185
rect 341 173 345 177
rect 533 194 537 198
rect 608 279 612 283
rect 751 279 755 283
rect 643 269 647 273
rect 584 251 588 255
rect 616 253 620 257
rect 653 253 657 257
rect 673 252 677 256
rect 728 271 732 275
rect 720 252 724 256
rect 644 236 648 240
rect 729 236 733 240
rect 806 272 811 276
rect 757 252 761 256
rect 840 279 844 283
rect 809 236 813 240
rect 848 254 852 258
rect 561 222 568 229
rect 645 206 650 211
rect 565 194 569 198
rect 636 194 640 198
rect 194 149 199 153
rect 214 148 219 153
rect 658 199 662 203
rect 677 184 681 188
rect 668 176 672 180
rect 721 199 725 203
rect 729 193 733 198
rect 658 168 662 172
rect 646 162 650 166
rect 728 158 733 165
rect -49 128 -45 132
rect -73 100 -69 104
rect -41 102 -37 106
rect -4 102 0 106
rect 16 101 20 105
rect 63 101 67 105
rect 94 128 98 132
rect 100 101 104 105
rect 77 85 81 89
rect 183 128 187 132
rect 152 85 156 89
rect 191 103 195 107
rect 194 75 202 82
rect 143 65 147 69
rect 20 33 24 37
rect 11 25 15 29
rect 138 46 144 52
rect 167 46 172 51
rect 192 46 197 51
rect 213 46 218 51
rect 280 130 284 134
rect 423 130 427 134
rect 316 111 320 115
rect 256 102 260 106
rect 288 104 292 108
rect 325 104 329 108
rect 345 103 349 107
rect 392 103 396 107
rect 316 87 320 91
rect 429 103 433 107
rect 512 130 516 134
rect 481 87 485 91
rect 520 105 524 109
rect 231 75 236 80
rect 521 76 525 80
rect 316 61 320 65
rect 316 43 320 47
rect 349 35 353 39
rect 340 27 344 31
rect 406 53 412 58
rect 494 53 499 58
rect 607 133 611 137
rect 750 133 754 137
rect 583 105 587 109
rect 615 107 619 111
rect 652 107 656 111
rect 672 106 676 110
rect 719 106 723 110
rect 756 106 760 110
rect 839 133 843 137
rect 808 90 812 94
rect 847 108 851 112
rect 561 76 565 80
rect 619 67 623 71
rect 558 53 563 58
rect 592 53 597 58
rect 389 20 394 25
rect 288 13 292 17
rect 676 38 680 42
rect 667 30 671 34
rect 724 55 730 60
rect 619 26 623 30
rect 288 -16 292 -12
rect 212 -52 217 -47
rect 260 -53 265 -48
rect 280 -64 284 -60
rect 390 -24 394 -19
rect 357 -36 361 -31
rect 353 -53 358 -48
rect 446 -36 450 -32
rect 438 -53 443 -48
rect 204 -75 211 -68
<< m3contact >>
rect 390 296 394 300
rect 409 275 413 279
<< psubstratepcontact >>
rect 36 363 40 367
rect 123 363 127 367
rect 216 363 220 367
rect 428 365 432 369
rect 521 365 525 369
rect 608 365 612 369
rect -70 224 -66 228
rect 8 224 12 228
rect 92 224 96 228
rect 162 224 166 228
rect 259 226 263 230
rect 337 226 341 230
rect 421 226 425 230
rect 491 226 495 230
rect 586 229 590 233
rect 664 229 668 233
rect 748 229 752 233
rect 818 229 822 233
rect 23 214 27 218
rect 51 214 55 218
rect 352 216 356 220
rect 380 216 384 220
rect 679 219 683 223
rect 707 219 711 223
rect -71 78 -67 82
rect 7 78 11 82
rect 91 78 95 82
rect 161 78 165 82
rect 258 80 262 84
rect 336 80 340 84
rect 420 80 424 84
rect 490 80 494 84
rect 585 83 589 87
rect 663 83 667 87
rect 747 83 751 87
rect 817 83 821 87
rect 22 68 26 72
rect 50 68 54 72
rect 351 70 355 74
rect 379 70 383 74
rect 678 73 682 77
rect 706 73 710 77
rect 223 -70 227 -66
rect 316 -70 320 -66
rect 403 -70 407 -66
<< nsubstratencontact >>
rect 36 303 40 307
rect 123 303 127 307
rect 216 303 220 307
rect 428 305 432 309
rect 521 305 525 309
rect 608 305 612 309
rect -70 284 -66 288
rect -56 284 -52 288
rect -42 284 -38 288
rect 41 284 45 288
rect 125 284 129 288
rect 162 284 166 288
rect 176 284 180 288
rect 190 284 194 288
rect 259 286 263 290
rect 273 286 277 290
rect 287 286 291 290
rect 370 286 374 290
rect 454 286 458 290
rect 491 286 495 290
rect 505 286 509 290
rect 519 286 523 290
rect 586 289 590 293
rect 600 289 604 293
rect 614 289 618 293
rect 697 289 701 293
rect 781 289 785 293
rect 818 289 822 293
rect 832 289 836 293
rect 846 289 850 293
rect 51 154 55 158
rect 380 156 384 160
rect 707 159 711 163
rect -71 138 -67 142
rect -57 138 -53 142
rect -43 138 -39 142
rect 40 138 44 142
rect 124 138 128 142
rect 161 138 165 142
rect 175 138 179 142
rect 189 138 193 142
rect 258 140 262 144
rect 272 140 276 144
rect 286 140 290 144
rect 369 140 373 144
rect 453 140 457 144
rect 490 140 494 144
rect 504 140 508 144
rect 518 140 522 144
rect 585 143 589 147
rect 599 143 603 147
rect 613 143 617 147
rect 696 143 700 147
rect 780 143 784 147
rect 817 143 821 147
rect 831 143 835 147
rect 845 143 849 147
rect 50 8 54 12
rect 379 10 383 14
rect 706 13 710 17
rect 223 -10 227 -6
rect 316 -10 320 -6
rect 403 -10 407 -6
<< psubstratepdiff >>
rect 427 369 433 370
rect 35 367 41 368
rect 35 363 36 367
rect 40 363 41 367
rect 35 362 41 363
rect 122 367 128 368
rect 122 363 123 367
rect 127 363 128 367
rect 122 362 128 363
rect 215 367 221 368
rect 215 363 216 367
rect 220 363 221 367
rect 427 365 428 369
rect 432 365 433 369
rect 427 364 433 365
rect 520 369 526 370
rect 520 365 521 369
rect 525 365 526 369
rect 215 362 221 363
rect 520 364 526 365
rect 607 369 613 370
rect 607 365 608 369
rect 612 365 613 369
rect 607 364 613 365
rect -71 228 -65 229
rect -71 224 -70 228
rect -66 224 -65 228
rect -71 223 -65 224
rect 7 228 13 229
rect 7 224 8 228
rect 12 224 13 228
rect 7 223 13 224
rect 91 228 97 229
rect 91 224 92 228
rect 96 224 97 228
rect 91 223 97 224
rect 258 230 264 231
rect 161 228 167 229
rect 161 224 162 228
rect 166 224 167 228
rect 161 223 167 224
rect 258 226 259 230
rect 263 226 264 230
rect 258 225 264 226
rect 336 230 342 231
rect 336 226 337 230
rect 341 226 342 230
rect 336 225 342 226
rect 420 230 426 231
rect 420 226 421 230
rect 425 226 426 230
rect 420 225 426 226
rect 585 233 591 234
rect 490 230 496 231
rect 490 226 491 230
rect 495 226 496 230
rect 490 225 496 226
rect 585 229 586 233
rect 590 229 591 233
rect 585 228 591 229
rect 663 233 669 234
rect 663 229 664 233
rect 668 229 669 233
rect 663 228 669 229
rect 747 233 753 234
rect 747 229 748 233
rect 752 229 753 233
rect 747 228 753 229
rect 817 233 823 234
rect 817 229 818 233
rect 822 229 823 233
rect 817 228 823 229
rect 678 223 712 224
rect 351 220 385 221
rect 22 218 56 219
rect 22 214 23 218
rect 27 214 51 218
rect 55 214 56 218
rect 351 216 352 220
rect 356 216 380 220
rect 384 216 385 220
rect 678 219 679 223
rect 683 219 707 223
rect 711 219 712 223
rect 678 218 712 219
rect 351 215 385 216
rect 22 213 56 214
rect -72 82 -66 83
rect -72 78 -71 82
rect -67 78 -66 82
rect -72 77 -66 78
rect 6 82 12 83
rect 6 78 7 82
rect 11 78 12 82
rect 6 77 12 78
rect 90 82 96 83
rect 90 78 91 82
rect 95 78 96 82
rect 90 77 96 78
rect 257 84 263 85
rect 160 82 166 83
rect 160 78 161 82
rect 165 78 166 82
rect 160 77 166 78
rect 257 80 258 84
rect 262 80 263 84
rect 257 79 263 80
rect 335 84 341 85
rect 335 80 336 84
rect 340 80 341 84
rect 335 79 341 80
rect 419 84 425 85
rect 419 80 420 84
rect 424 80 425 84
rect 419 79 425 80
rect 584 87 590 88
rect 489 84 495 85
rect 489 80 490 84
rect 494 80 495 84
rect 489 79 495 80
rect 584 83 585 87
rect 589 83 590 87
rect 584 82 590 83
rect 662 87 668 88
rect 662 83 663 87
rect 667 83 668 87
rect 662 82 668 83
rect 746 87 752 88
rect 746 83 747 87
rect 751 83 752 87
rect 746 82 752 83
rect 816 87 822 88
rect 816 83 817 87
rect 821 83 822 87
rect 816 82 822 83
rect 677 77 711 78
rect 350 74 384 75
rect 21 72 55 73
rect 21 68 22 72
rect 26 68 50 72
rect 54 68 55 72
rect 350 70 351 74
rect 355 70 379 74
rect 383 70 384 74
rect 677 73 678 77
rect 682 73 706 77
rect 710 73 711 77
rect 677 72 711 73
rect 350 69 384 70
rect 21 67 55 68
rect 222 -66 228 -65
rect 222 -70 223 -66
rect 227 -70 228 -66
rect 222 -71 228 -70
rect 315 -66 321 -65
rect 315 -70 316 -66
rect 320 -70 321 -66
rect 315 -71 321 -70
rect 402 -66 408 -65
rect 402 -70 403 -66
rect 407 -70 408 -66
rect 402 -71 408 -70
<< nsubstratendiff >>
rect 35 307 41 308
rect 122 307 128 308
rect 427 309 433 310
rect 520 309 526 310
rect 607 309 613 310
rect 215 307 221 308
rect 35 303 36 307
rect 40 303 41 307
rect 35 302 41 303
rect 122 303 123 307
rect 127 303 128 307
rect 122 302 128 303
rect 215 303 216 307
rect 220 303 221 307
rect 427 305 428 309
rect 432 305 433 309
rect 427 304 433 305
rect 520 305 521 309
rect 525 305 526 309
rect 520 304 526 305
rect 607 305 608 309
rect 612 305 613 309
rect 607 304 613 305
rect 215 302 221 303
rect 258 290 292 291
rect -71 288 -37 289
rect -71 284 -70 288
rect -66 284 -56 288
rect -52 284 -42 288
rect -38 284 -37 288
rect 40 288 46 289
rect -71 283 -37 284
rect 40 284 41 288
rect 45 284 46 288
rect 124 288 130 289
rect 40 283 46 284
rect 124 284 125 288
rect 129 284 130 288
rect 161 288 195 289
rect 124 283 130 284
rect 161 284 162 288
rect 166 284 176 288
rect 180 284 190 288
rect 194 284 195 288
rect 258 286 259 290
rect 263 286 273 290
rect 277 286 287 290
rect 291 286 292 290
rect 369 290 375 291
rect 258 285 292 286
rect 161 283 195 284
rect 369 286 370 290
rect 374 286 375 290
rect 453 290 459 291
rect 369 285 375 286
rect 453 286 454 290
rect 458 286 459 290
rect 490 290 524 291
rect 453 285 459 286
rect 490 286 491 290
rect 495 286 505 290
rect 509 286 519 290
rect 523 286 524 290
rect 585 289 586 293
rect 590 289 600 293
rect 604 289 614 293
rect 618 289 619 293
rect 696 293 702 294
rect 585 288 619 289
rect 490 285 524 286
rect 696 289 697 293
rect 701 289 702 293
rect 780 293 786 294
rect 696 288 702 289
rect 780 289 781 293
rect 785 289 786 293
rect 817 293 851 294
rect 780 288 786 289
rect 817 289 818 293
rect 822 289 832 293
rect 836 289 846 293
rect 850 289 851 293
rect 817 288 851 289
rect 50 158 56 159
rect 706 163 712 164
rect 379 160 385 161
rect 50 154 51 158
rect 55 154 56 158
rect 379 156 380 160
rect 384 156 385 160
rect 706 159 707 163
rect 711 159 712 163
rect 706 158 712 159
rect 379 155 385 156
rect 50 153 56 154
rect 584 147 618 148
rect 257 144 291 145
rect -72 142 -38 143
rect -72 138 -71 142
rect -67 138 -57 142
rect -53 138 -43 142
rect -39 138 -38 142
rect 39 142 45 143
rect -72 137 -38 138
rect 39 138 40 142
rect 44 138 45 142
rect 123 142 129 143
rect 39 137 45 138
rect 123 138 124 142
rect 128 138 129 142
rect 160 142 194 143
rect 123 137 129 138
rect 160 138 161 142
rect 165 138 175 142
rect 179 138 189 142
rect 193 138 194 142
rect 257 140 258 144
rect 262 140 272 144
rect 276 140 286 144
rect 290 140 291 144
rect 368 144 374 145
rect 257 139 291 140
rect 160 137 194 138
rect 368 140 369 144
rect 373 140 374 144
rect 452 144 458 145
rect 368 139 374 140
rect 452 140 453 144
rect 457 140 458 144
rect 489 144 523 145
rect 452 139 458 140
rect 489 140 490 144
rect 494 140 504 144
rect 508 140 518 144
rect 522 140 523 144
rect 584 143 585 147
rect 589 143 599 147
rect 603 143 613 147
rect 617 143 618 147
rect 695 147 701 148
rect 584 142 618 143
rect 489 139 523 140
rect 695 143 696 147
rect 700 143 701 147
rect 779 147 785 148
rect 695 142 701 143
rect 779 143 780 147
rect 784 143 785 147
rect 816 147 850 148
rect 779 142 785 143
rect 816 143 817 147
rect 821 143 831 147
rect 835 143 845 147
rect 849 143 850 147
rect 816 142 850 143
rect 49 12 55 13
rect 705 17 711 18
rect 378 14 384 15
rect 49 8 50 12
rect 54 8 55 12
rect 378 10 379 14
rect 383 10 384 14
rect 705 13 706 17
rect 710 13 711 17
rect 705 12 711 13
rect 378 9 384 10
rect 49 7 55 8
rect 222 -6 228 -5
rect 222 -10 223 -6
rect 227 -10 228 -6
rect 315 -6 321 -5
rect 315 -10 316 -6
rect 320 -10 321 -6
rect 402 -6 408 -5
rect 402 -10 403 -6
rect 407 -10 408 -6
rect 222 -11 228 -10
rect 315 -11 321 -10
rect 402 -11 408 -10
<< pad >>
rect 63 297 67 301
<< labels >>
rlabel metal1 368 220 368 220 2 vss
rlabel metal1 602 229 602 229 6 vss
rlabel metal1 834 293 834 293 6 vdd
rlabel metal1 695 223 695 223 2 vss
rlabel metal1 695 159 695 159 2 vdd
rlabel metal1 694 13 694 13 2 vdd
rlabel metal1 694 77 694 77 2 vss
rlabel metal1 833 83 833 83 6 vss
rlabel metal1 833 147 833 147 6 vdd
rlabel metal1 601 147 601 147 6 vdd
rlabel metal1 601 83 601 83 6 vss
rlabel metal1 691 147 691 147 6 vdd
rlabel metal1 367 74 367 74 2 vss
rlabel metal1 506 80 506 80 6 vss
rlabel metal1 506 144 506 144 6 vdd
rlabel metal1 274 144 274 144 6 vdd
rlabel metal1 274 80 274 80 6 vss
rlabel metal1 448 144 448 144 6 vdd
rlabel metal1 448 80 448 80 6 vss
rlabel metal1 38 8 38 8 2 vdd
rlabel metal1 -55 142 -55 142 6 vdd
rlabel metal1 -55 78 -55 78 6 vss
rlabel metal1 119 142 119 142 6 vdd
rlabel metal1 119 78 119 78 6 vss
rlabel m2contact 4 347 4 347 1 q0_M2
rlabel metal1 32 343 32 343 1 q0b2_n_M2
rlabel metal1 40 339 40 339 1 q0b2_M2
rlabel metal1 119 344 119 344 1 q0b1_n_M2
rlabel metal1 127 343 127 343 1 q0b1_M2
rlabel metal1 212 346 212 346 1 q0b0_n_M2
rlabel metal1 219 345 219 345 1 a0_M2
rlabel metal1 332 352 332 352 1 b2_M2
rlabel metal1 333 312 333 312 1 b0_M2
rlabel metal1 333 331 333 331 1 b1_M2
rlabel metal1 529 357 529 357 1 q1b1_M2
rlabel metal1 607 346 607 346 1 q1b2_M2
rlabel metal1 616 346 616 346 1 q1b2_n_M2
rlabel m2contact 643 349 643 349 1 q1_M2
rlabel metal1 832 257 832 257 1 zc1_n_3_M2
rlabel metal1 818 257 818 257 1 c1_3_M2
rlabel metal1 804 261 804 261 1 s_fa3_M2
rlabel ntransistor 797 244 797 244 1 s_fa3_n_M2
rlabel metal1 720 261 720 261 1 so_3_M2
rlabel metal1 607 261 607 261 1 co_n3_M2
rlabel metal1 594 241 594 241 1 co_3_M2
rlabel metal1 505 254 505 254 1 zc1_2_n_M2
rlabel metal1 491 254 491 254 1 c1_2_M2
rlabel pdcontact 467 271 467 271 1 s_fa2_M2
rlabel metal1 455 254 455 254 1 cn2_M2
rlabel ntransistor 470 241 470 241 1 son_2_M2
rlabel metal1 393 258 393 258 1 so_2_M2
rlabel polycontact 376 255 376 255 1 bn_2_M2
rlabel polycontact 385 255 385 255 1 an_2_M2
rlabel metal1 280 257 280 257 1 co_n2_M2
rlabel metal1 267 238 267 238 1 co_2_M2
rlabel metal1 176 252 176 252 1 zc1_n1_M2
rlabel metal1 162 252 162 252 1 c1_1_M2
rlabel metal1 148 256 148 256 1 a1_M2
rlabel ntransistor 141 239 141 239 1 a1_1_M2
rlabel metal1 64 256 64 256 1 so_1_M2
rlabel ntransistor 57 240 57 240 1 an_1_M2
rlabel metal1 52 277 52 277 1 bn_1_M1
rlabel metal1 -62 236 -62 236 1 co_1_M2
rlabel metal1 -49 256 -49 256 1 co_n1_M2
rlabel metal1 47 184 47 184 1 c_fa1_n_M2
rlabel metal1 55 184 55 184 1 c_fa1_M2
rlabel metal1 376 188 376 188 1 c_fa2_n_M2
rlabel metal1 384 192 384 192 1 c_fa2_M2
rlabel metal1 703 191 703 191 1 c_fa3_n_M2
rlabel metal1 711 195 711 195 1 c_fa3_M2
rlabel metal1 831 111 831 111 1 zc1_6_n_M2
rlabel metal1 817 111 817 111 1 c1_6_M2
rlabel ntransistor 796 98 796 98 1 s_fa_6_n_M2
rlabel metal1 803 115 803 115 1 a2_M2
rlabel metal1 779 132 779 132 1 cn_6_M2
rlabel metal1 719 115 719 115 1 so_6_M2
rlabel ptransistor 703 120 703 120 1 an_6_M2
rlabel metal1 664 109 664 109 1 bn_6_M2
rlabel metal1 606 115 606 115 1 co_n_6_M2
rlabel metal1 593 95 593 95 1 co_6_M2
rlabel metal1 504 108 504 108 1 zc1_n_5_M2
rlabel metal1 490 108 490 108 1 c1_5_M2
rlabel ntransistor 469 95 469 95 1 s_fa_5_n_M2
rlabel metal1 476 112 476 112 1 a3_M2
rlabel metal1 452 128 452 128 1 cn_5_M2
rlabel metal1 380 133 380 133 1 bn_5_M2
rlabel ptransistor 376 117 376 117 1 an_5_M2
rlabel metal1 392 112 392 112 1 so_5_M2
rlabel metal1 175 106 175 106 1 zc1_4_M2
rlabel metal1 161 106 161 106 1 c1_4_M2
rlabel metal1 147 110 147 110 1 a4_M2
rlabel ntransistor 140 93 140 93 1 s_fa4_n_M2
rlabel metal1 123 126 123 126 1 cn_1_M2
rlabel metal1 40 125 40 125 1 bn4_M2
rlabel ptransistor 47 115 47 115 1 an4_M2
rlabel metal1 63 110 63 110 1 so_4_M2
rlabel metal1 -50 110 -50 110 1 co_n4_M2
rlabel metal1 -63 90 -63 90 1 co_4_M2
rlabel polycontact 46 43 46 43 1 a5_n_M2
rlabel metal1 54 44 54 44 1 a5_M2
rlabel metal1 375 42 375 42 1 c_fa5_n_M2
rlabel metal1 383 46 383 46 1 c_fa5_M2
rlabel metal1 702 45 702 45 1 c_fa6_n_M2
rlabel metal1 710 49 710 49 1 c_fa6_M2
rlabel metal1 245 -59 245 -59 1 q2b2_n_M2
rlabel metal1 223 -60 223 -60 1 q2b2_M2
rlabel metal1 315 -48 315 -48 1 q2b1_M2
rlabel metal1 324 -48 324 -48 1 q2b1_n_M2
rlabel m2contact 440 -50 440 -50 1 q2_M2
rlabel metal1 412 -49 412 -49 1 q2b0_n_M2
rlabel metal1 403 -48 403 -48 1 q2b0_M2
rlabel metal1 427 350 427 350 1 q1b0_M2
rlabel metal1 436 336 436 336 1 q1b0_n_M2
rlabel metal1 781 279 781 279 1 cn_3_M2
rlabel ptransistor 704 266 704 266 1 an3_M2
rlabel metal1 708 282 708 282 1 bn3_M2
rlabel metal1 279 112 279 112 1 co_5_M2
rlabel metal1 529 335 529 335 1 q1b1_n_M2
rlabel metal1 -96 342 -96 342 1 q0_M2
rlabel metal2 -98 390 -98 390 5 q1_M2
rlabel metal2 207 397 207 397 1 b0_M2
rlabel metal2 206 404 206 404 1 b1_M2
rlabel metal2 209 411 209 411 5 b2_M2
rlabel metal1 183 -50 184 -50 1 q2_M2
<< end >>
