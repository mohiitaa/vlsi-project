magic
tech scmos
timestamp 1521735912
<< pwell >>
rect 174 71 317 102
rect 148 66 317 71
rect 329 66 447 102
rect 148 39 250 66
rect 260 40 308 66
<< nwell >>
rect 174 102 317 146
rect 329 102 447 146
rect 148 38 250 39
rect 260 38 308 40
rect 148 -4 308 38
rect 148 -5 261 -4
<< polysilicon >>
rect 266 136 268 140
rect 190 128 196 129
rect 180 120 182 125
rect 190 124 191 128
rect 195 124 196 128
rect 190 123 196 124
rect 190 118 192 123
rect 200 118 202 123
rect 251 120 257 121
rect 251 116 252 120
rect 256 116 257 120
rect 251 115 257 116
rect 180 105 182 108
rect 190 105 192 108
rect 180 104 186 105
rect 180 100 181 104
rect 185 100 186 104
rect 190 102 194 105
rect 180 99 186 100
rect 180 91 182 99
rect 192 88 194 102
rect 200 97 202 108
rect 255 106 257 115
rect 302 136 304 140
rect 350 136 352 140
rect 282 127 284 131
rect 292 127 294 131
rect 335 120 341 121
rect 335 116 336 120
rect 340 116 341 120
rect 335 115 341 116
rect 266 106 268 109
rect 282 106 284 109
rect 292 106 294 109
rect 302 106 304 109
rect 255 104 268 106
rect 274 104 284 106
rect 288 105 294 106
rect 199 96 205 97
rect 258 96 260 104
rect 274 100 276 104
rect 288 101 289 105
rect 293 101 294 105
rect 288 100 294 101
rect 298 105 304 106
rect 298 101 299 105
rect 303 101 304 105
rect 339 106 341 115
rect 386 136 388 140
rect 366 127 368 131
rect 376 127 378 131
rect 422 128 428 129
rect 412 120 414 125
rect 422 124 423 128
rect 427 124 428 128
rect 422 123 428 124
rect 350 106 352 109
rect 366 106 368 109
rect 376 106 378 109
rect 386 106 388 109
rect 422 118 424 123
rect 432 118 434 123
rect 339 104 352 106
rect 358 104 368 106
rect 372 105 378 106
rect 298 100 304 101
rect 267 99 276 100
rect 199 92 200 96
rect 204 92 205 96
rect 199 91 205 92
rect 199 88 201 91
rect 180 81 182 85
rect 267 95 268 99
rect 272 95 276 99
rect 292 96 294 100
rect 267 94 276 95
rect 274 91 276 94
rect 284 91 286 96
rect 292 94 296 96
rect 294 91 296 94
rect 301 91 303 100
rect 342 96 344 104
rect 358 100 360 104
rect 372 101 373 105
rect 377 101 378 105
rect 372 100 378 101
rect 382 105 388 106
rect 382 101 383 105
rect 387 101 388 105
rect 382 100 388 101
rect 412 105 414 108
rect 422 105 424 108
rect 412 104 418 105
rect 412 100 413 104
rect 417 100 418 104
rect 422 102 426 105
rect 351 99 360 100
rect 258 84 260 87
rect 258 82 263 84
rect 192 74 194 79
rect 199 74 201 79
rect 261 74 263 82
rect 274 78 276 82
rect 284 74 286 82
rect 351 95 352 99
rect 356 95 360 99
rect 376 96 378 100
rect 351 94 360 95
rect 358 91 360 94
rect 368 91 370 96
rect 376 94 380 96
rect 378 91 380 94
rect 385 91 387 100
rect 412 99 418 100
rect 412 91 414 99
rect 342 84 344 87
rect 342 82 347 84
rect 294 74 296 79
rect 301 74 303 79
rect 261 72 286 74
rect 345 74 347 82
rect 358 78 360 82
rect 368 74 370 82
rect 424 88 426 102
rect 432 97 434 108
rect 431 96 437 97
rect 431 92 432 96
rect 436 92 437 96
rect 431 91 437 92
rect 431 88 433 91
rect 412 81 414 85
rect 378 74 380 79
rect 385 74 387 79
rect 345 72 370 74
rect 424 74 426 79
rect 431 74 433 79
rect 169 65 171 69
rect 180 65 182 69
rect 187 65 189 69
rect 169 42 171 51
rect 207 59 209 64
rect 217 59 219 64
rect 227 62 229 67
rect 237 65 239 69
rect 273 57 275 61
rect 283 57 285 61
rect 293 57 295 61
rect 180 42 182 45
rect 187 42 189 45
rect 207 42 209 45
rect 217 42 219 45
rect 167 41 173 42
rect 167 37 168 41
rect 172 37 173 41
rect 167 36 173 37
rect 177 41 183 42
rect 177 37 178 41
rect 182 37 183 41
rect 177 36 183 37
rect 187 41 209 42
rect 187 37 188 41
rect 192 37 195 41
rect 199 37 209 41
rect 187 36 209 37
rect 213 41 219 42
rect 213 37 214 41
rect 218 37 219 41
rect 213 36 219 37
rect 227 39 229 52
rect 237 49 239 52
rect 233 48 239 49
rect 233 44 234 48
rect 238 44 239 48
rect 233 43 239 44
rect 273 43 275 51
rect 227 38 233 39
rect 169 33 171 36
rect 179 33 181 36
rect 189 33 191 36
rect 207 33 209 36
rect 214 33 216 36
rect 227 35 228 38
rect 224 34 228 35
rect 232 34 233 38
rect 224 33 233 34
rect 224 30 226 33
rect 237 30 239 43
rect 269 42 275 43
rect 283 42 285 51
rect 293 42 295 51
rect 269 38 270 42
rect 274 38 275 42
rect 289 41 295 42
rect 269 37 275 38
rect 224 12 226 17
rect 169 1 171 5
rect 179 1 181 5
rect 189 1 191 5
rect 207 3 209 8
rect 214 3 216 8
rect 273 24 275 37
rect 283 35 285 38
rect 289 37 290 41
rect 294 37 295 41
rect 289 36 295 37
rect 279 34 285 35
rect 279 30 280 34
rect 284 30 285 34
rect 279 29 285 30
rect 280 24 282 29
rect 293 27 295 36
rect 293 11 295 15
rect 237 1 239 5
rect 273 2 275 6
rect 280 2 282 6
<< ndiffusion >>
rect 173 90 180 91
rect 173 86 174 90
rect 178 86 180 90
rect 173 85 180 86
rect 182 88 190 91
rect 251 95 258 96
rect 251 91 252 95
rect 256 91 258 95
rect 251 90 258 91
rect 182 85 192 88
rect 184 79 192 85
rect 194 79 199 88
rect 201 87 208 88
rect 253 87 258 90
rect 260 91 265 96
rect 335 95 342 96
rect 335 91 336 95
rect 340 91 342 95
rect 260 87 274 91
rect 201 83 203 87
rect 207 83 208 87
rect 201 82 208 83
rect 265 83 266 87
rect 270 83 274 87
rect 265 82 274 83
rect 276 90 284 91
rect 276 86 278 90
rect 282 86 284 90
rect 276 82 284 86
rect 286 88 294 91
rect 286 84 288 88
rect 292 84 294 88
rect 286 82 294 84
rect 201 79 206 82
rect 184 78 190 79
rect 184 74 185 78
rect 189 74 190 78
rect 184 73 190 74
rect 289 79 294 82
rect 296 79 301 91
rect 303 79 311 91
rect 335 90 342 91
rect 337 87 342 90
rect 344 91 349 96
rect 344 87 358 91
rect 349 83 350 87
rect 354 83 358 87
rect 349 82 358 83
rect 360 90 368 91
rect 360 86 362 90
rect 366 86 368 90
rect 360 82 368 86
rect 370 88 378 91
rect 370 84 372 88
rect 376 84 378 88
rect 370 82 378 84
rect 305 78 311 79
rect 305 74 306 78
rect 310 74 311 78
rect 305 73 311 74
rect 373 79 378 82
rect 380 79 385 91
rect 387 79 395 91
rect 405 90 412 91
rect 405 86 406 90
rect 410 86 412 90
rect 405 85 412 86
rect 414 88 422 91
rect 414 85 424 88
rect 416 79 424 85
rect 426 79 431 88
rect 433 87 440 88
rect 433 83 435 87
rect 439 83 440 87
rect 433 82 440 83
rect 433 79 438 82
rect 389 78 395 79
rect 389 74 390 78
rect 394 74 395 78
rect 389 73 395 74
rect 416 78 422 79
rect 416 74 417 78
rect 421 74 422 78
rect 416 73 422 74
rect 164 58 169 65
rect 162 57 169 58
rect 162 53 163 57
rect 167 53 169 57
rect 162 51 169 53
rect 171 64 180 65
rect 171 60 174 64
rect 178 60 180 64
rect 171 51 180 60
rect 173 45 180 51
rect 182 45 187 65
rect 189 58 194 65
rect 232 62 237 65
rect 222 59 227 62
rect 189 57 196 58
rect 189 53 191 57
rect 195 53 196 57
rect 189 52 196 53
rect 200 57 207 59
rect 200 53 201 57
rect 205 53 207 57
rect 189 45 194 52
rect 200 50 207 53
rect 200 46 201 50
rect 205 46 207 50
rect 200 45 207 46
rect 209 50 217 59
rect 209 46 211 50
rect 215 46 217 50
rect 209 45 217 46
rect 219 58 227 59
rect 219 54 221 58
rect 225 54 227 58
rect 219 52 227 54
rect 229 61 237 62
rect 229 57 231 61
rect 235 57 237 61
rect 229 52 237 57
rect 239 58 244 65
rect 239 57 246 58
rect 239 53 241 57
rect 245 53 246 57
rect 239 52 246 53
rect 266 56 273 57
rect 266 52 267 56
rect 271 52 273 56
rect 219 45 224 52
rect 266 51 273 52
rect 275 56 283 57
rect 275 52 277 56
rect 281 52 283 56
rect 275 51 283 52
rect 285 56 293 57
rect 285 52 287 56
rect 291 52 293 56
rect 285 51 293 52
rect 295 56 302 57
rect 295 52 297 56
rect 301 52 302 56
rect 295 51 302 52
<< pdiffusion >>
rect 175 114 180 120
rect 173 113 180 114
rect 173 109 174 113
rect 178 109 180 113
rect 173 108 180 109
rect 182 118 188 120
rect 182 113 190 118
rect 182 109 184 113
rect 188 109 190 113
rect 182 108 190 109
rect 192 113 200 118
rect 192 109 194 113
rect 198 109 200 113
rect 192 108 200 109
rect 202 117 209 118
rect 202 113 204 117
rect 208 113 209 117
rect 261 115 266 136
rect 202 108 209 113
rect 259 114 266 115
rect 259 110 260 114
rect 264 110 266 114
rect 259 109 266 110
rect 268 135 280 136
rect 268 131 270 135
rect 274 131 280 135
rect 268 128 280 131
rect 268 124 270 128
rect 274 127 280 128
rect 297 127 302 136
rect 274 124 282 127
rect 268 109 282 124
rect 284 114 292 127
rect 284 110 286 114
rect 290 110 292 114
rect 284 109 292 110
rect 294 121 302 127
rect 294 117 296 121
rect 300 117 302 121
rect 294 109 302 117
rect 304 130 309 136
rect 304 129 311 130
rect 304 125 306 129
rect 310 125 311 129
rect 304 124 311 125
rect 304 109 309 124
rect 345 115 350 136
rect 343 114 350 115
rect 343 110 344 114
rect 348 110 350 114
rect 343 109 350 110
rect 352 135 364 136
rect 352 131 354 135
rect 358 131 364 135
rect 352 128 364 131
rect 352 124 354 128
rect 358 127 364 128
rect 381 127 386 136
rect 358 124 366 127
rect 352 109 366 124
rect 368 114 376 127
rect 368 110 370 114
rect 374 110 376 114
rect 368 109 376 110
rect 378 121 386 127
rect 378 117 380 121
rect 384 117 386 121
rect 378 109 386 117
rect 388 130 393 136
rect 388 129 395 130
rect 388 125 390 129
rect 394 125 395 129
rect 388 124 395 125
rect 388 109 393 124
rect 407 114 412 120
rect 405 113 412 114
rect 405 109 406 113
rect 410 109 412 113
rect 405 108 412 109
rect 414 118 420 120
rect 414 113 422 118
rect 414 109 416 113
rect 420 109 422 113
rect 414 108 422 109
rect 424 113 432 118
rect 424 109 426 113
rect 430 109 432 113
rect 424 108 432 109
rect 434 117 441 118
rect 434 113 436 117
rect 440 113 441 117
rect 434 108 441 113
rect 162 32 169 33
rect 162 28 163 32
rect 167 28 169 32
rect 162 25 169 28
rect 162 21 163 25
rect 167 21 169 25
rect 162 20 169 21
rect 164 5 169 20
rect 171 17 179 33
rect 171 13 173 17
rect 177 13 179 17
rect 171 10 179 13
rect 171 6 173 10
rect 177 6 179 10
rect 171 5 179 6
rect 181 25 189 33
rect 181 21 183 25
rect 187 21 189 25
rect 181 18 189 21
rect 181 14 183 18
rect 187 14 189 18
rect 181 5 189 14
rect 191 17 207 33
rect 191 13 195 17
rect 199 13 207 17
rect 191 10 207 13
rect 191 6 195 10
rect 199 8 207 10
rect 209 8 214 33
rect 216 30 221 33
rect 216 29 224 30
rect 216 25 218 29
rect 222 25 224 29
rect 216 17 224 25
rect 226 17 237 30
rect 216 8 221 17
rect 228 10 237 17
rect 199 6 205 8
rect 191 5 205 6
rect 228 6 230 10
rect 234 6 237 10
rect 228 5 237 6
rect 239 29 246 30
rect 239 25 241 29
rect 245 25 246 29
rect 239 22 246 25
rect 285 24 293 27
rect 239 18 241 22
rect 245 18 246 22
rect 268 19 273 24
rect 239 17 246 18
rect 266 18 273 19
rect 239 5 244 17
rect 266 14 267 18
rect 271 14 273 18
rect 266 13 273 14
rect 268 6 273 13
rect 275 6 280 24
rect 282 15 293 24
rect 295 21 300 27
rect 295 20 302 21
rect 295 16 297 20
rect 301 16 302 20
rect 295 15 302 16
rect 282 11 291 15
rect 282 7 285 11
rect 289 7 291 11
rect 282 6 291 7
<< metal1 >>
rect 139 138 445 142
rect 139 134 175 138
rect 179 134 189 138
rect 193 134 203 138
rect 207 135 286 138
rect 207 134 270 135
rect 139 23 143 134
rect 173 114 177 121
rect 173 113 178 114
rect 173 109 174 113
rect 181 113 185 134
rect 188 128 201 129
rect 188 124 191 128
rect 195 124 197 128
rect 188 123 201 124
rect 188 116 194 123
rect 204 117 208 134
rect 274 134 286 135
rect 290 135 370 138
rect 290 134 354 135
rect 251 123 263 129
rect 270 128 274 131
rect 358 134 370 135
rect 374 134 407 138
rect 411 134 421 138
rect 425 134 435 138
rect 439 134 445 138
rect 284 125 306 129
rect 310 125 311 129
rect 335 128 347 129
rect 284 124 288 125
rect 270 123 274 124
rect 251 120 256 123
rect 251 119 252 120
rect 181 109 184 113
rect 188 109 189 113
rect 193 109 194 113
rect 198 109 199 113
rect 204 112 208 113
rect 243 116 252 119
rect 277 120 288 124
rect 335 124 340 128
rect 344 124 347 128
rect 335 123 347 124
rect 354 128 358 131
rect 368 125 390 129
rect 394 125 395 129
rect 368 124 372 125
rect 354 123 358 124
rect 277 116 281 120
rect 295 117 296 121
rect 300 117 311 121
rect 173 108 178 109
rect 173 100 177 108
rect 193 104 199 109
rect 180 100 181 104
rect 185 100 199 104
rect 205 102 209 105
rect 243 102 246 116
rect 251 115 256 116
rect 260 114 281 116
rect 173 91 177 96
rect 173 90 178 91
rect 173 86 174 90
rect 178 86 185 89
rect 173 83 185 86
rect 189 87 193 100
rect 252 110 260 111
rect 264 112 281 114
rect 252 107 264 110
rect 205 96 209 98
rect 196 92 200 96
rect 204 92 209 96
rect 196 91 209 92
rect 252 95 256 107
rect 277 105 281 112
rect 285 110 286 114
rect 290 113 291 114
rect 290 110 302 113
rect 285 109 302 110
rect 298 106 302 109
rect 298 105 303 106
rect 266 99 272 104
rect 277 101 289 105
rect 293 101 294 105
rect 298 101 299 105
rect 266 97 268 99
rect 259 95 268 97
rect 298 100 303 101
rect 307 101 311 117
rect 335 120 340 123
rect 335 116 336 120
rect 361 120 372 124
rect 361 116 365 120
rect 379 117 380 121
rect 384 117 395 121
rect 335 115 340 116
rect 344 114 365 116
rect 336 110 344 111
rect 348 112 365 114
rect 336 107 348 110
rect 298 96 302 100
rect 259 91 272 95
rect 278 92 302 96
rect 307 97 309 101
rect 252 90 256 91
rect 278 90 282 92
rect 189 83 203 87
rect 207 83 208 87
rect 265 83 266 87
rect 270 83 271 87
rect 307 88 311 97
rect 336 95 340 107
rect 361 105 365 112
rect 369 110 370 114
rect 374 113 375 114
rect 374 110 386 113
rect 369 109 386 110
rect 382 106 386 109
rect 382 105 387 106
rect 350 99 356 104
rect 361 101 373 105
rect 377 101 378 105
rect 382 101 383 105
rect 350 97 352 99
rect 343 95 352 97
rect 382 100 387 101
rect 382 96 386 100
rect 343 91 356 95
rect 362 92 386 96
rect 336 90 340 91
rect 362 90 366 92
rect 278 85 282 86
rect 287 84 288 88
rect 292 84 311 88
rect 265 78 271 83
rect 349 83 350 87
rect 354 83 355 87
rect 391 88 395 117
rect 405 114 409 121
rect 405 113 410 114
rect 405 109 406 113
rect 413 113 417 134
rect 420 128 433 129
rect 420 124 423 128
rect 427 124 429 128
rect 420 123 433 124
rect 420 116 426 123
rect 436 117 440 134
rect 413 109 416 113
rect 420 109 421 113
rect 425 109 426 113
rect 430 109 431 113
rect 436 112 440 113
rect 405 108 410 109
rect 405 100 409 108
rect 425 104 431 109
rect 412 100 413 104
rect 417 100 431 104
rect 437 103 441 105
rect 362 85 366 86
rect 371 84 372 88
rect 376 84 395 88
rect 399 97 409 100
rect 399 85 402 97
rect 349 78 355 83
rect 405 91 409 97
rect 405 90 410 91
rect 405 86 406 90
rect 410 86 417 89
rect 405 83 417 86
rect 421 87 425 100
rect 437 96 441 99
rect 428 92 432 96
rect 436 92 441 96
rect 428 91 441 92
rect 421 83 435 87
rect 439 83 440 87
rect 172 74 175 78
rect 179 74 185 78
rect 189 74 253 78
rect 257 74 306 78
rect 310 74 337 78
rect 341 74 390 78
rect 394 74 407 78
rect 411 74 417 78
rect 421 74 445 78
rect 172 71 445 74
rect 150 70 445 71
rect 150 64 250 70
rect 262 68 306 70
rect 262 64 268 68
rect 272 64 296 68
rect 300 64 306 68
rect 150 63 174 64
rect 173 60 174 63
rect 178 63 250 64
rect 178 60 179 63
rect 231 61 235 63
rect 201 57 221 58
rect 138 3 143 23
rect 161 53 163 57
rect 167 53 183 57
rect 186 53 191 57
rect 195 53 196 57
rect 205 54 221 57
rect 225 54 226 58
rect 231 56 235 57
rect 241 57 246 58
rect 161 33 165 53
rect 186 49 190 53
rect 201 50 205 53
rect 245 53 246 57
rect 241 52 246 53
rect 266 56 272 64
rect 266 52 267 56
rect 271 52 272 56
rect 277 56 281 57
rect 286 56 292 64
rect 286 52 287 56
rect 291 52 292 56
rect 297 56 302 59
rect 301 52 302 56
rect 170 45 190 49
rect 170 42 174 45
rect 168 41 174 42
rect 172 37 174 41
rect 168 36 174 37
rect 161 32 167 33
rect 161 28 163 32
rect 161 25 167 28
rect 161 21 163 25
rect 170 25 174 36
rect 178 41 182 42
rect 194 41 198 50
rect 210 46 211 50
rect 215 48 225 50
rect 215 46 234 48
rect 201 45 205 46
rect 221 44 234 46
rect 238 44 239 48
rect 210 41 218 42
rect 185 37 188 41
rect 192 37 195 41
rect 199 37 200 41
rect 210 37 214 41
rect 178 33 182 37
rect 210 36 218 37
rect 210 33 215 36
rect 221 33 225 44
rect 177 29 215 33
rect 218 29 225 33
rect 228 38 232 39
rect 228 25 232 34
rect 242 30 246 52
rect 277 49 281 52
rect 297 51 302 52
rect 277 45 294 49
rect 170 21 183 25
rect 187 21 210 25
rect 218 24 222 25
rect 226 21 232 25
rect 241 29 246 30
rect 266 33 270 43
rect 274 38 279 42
rect 290 41 294 45
rect 274 30 280 34
rect 284 30 287 34
rect 245 25 246 29
rect 241 22 246 25
rect 161 20 167 21
rect 183 18 187 21
rect 172 13 173 17
rect 177 13 178 17
rect 206 17 230 21
rect 245 18 246 22
rect 274 24 278 30
rect 290 26 294 37
rect 261 21 278 24
rect 282 22 294 26
rect 282 18 286 22
rect 298 21 302 51
rect 297 20 302 21
rect 241 17 246 18
rect 183 13 187 14
rect 194 13 195 17
rect 199 13 200 17
rect 233 13 246 17
rect 266 14 267 18
rect 271 14 286 18
rect 289 16 297 18
rect 301 16 302 20
rect 289 14 302 16
rect 172 10 178 13
rect 172 7 173 10
rect 150 6 173 7
rect 177 7 178 10
rect 194 10 200 13
rect 194 7 195 10
rect 177 6 195 7
rect 199 7 200 10
rect 229 7 230 10
rect 199 6 230 7
rect 234 7 235 10
rect 284 8 285 11
rect 262 7 285 8
rect 289 8 290 11
rect 289 7 296 8
rect 234 6 250 7
rect 150 3 250 6
rect 262 4 296 7
rect 300 4 306 8
rect 262 3 306 4
rect 138 0 306 3
rect 138 -1 262 0
<< metal2 >>
rect 201 125 266 128
rect 166 97 173 100
rect 166 32 169 97
rect 209 98 242 101
rect 262 101 265 125
rect 334 124 340 127
rect 344 125 429 128
rect 334 100 337 124
rect 313 97 346 100
rect 326 93 329 97
rect 334 93 337 97
rect 438 93 441 99
rect 326 90 441 93
rect 334 56 337 90
rect 402 81 403 84
rect 179 53 337 56
rect 400 33 403 81
rect 166 29 260 32
rect 270 30 413 33
rect 257 25 260 29
<< ntransistor >>
rect 180 85 182 91
rect 192 79 194 88
rect 199 79 201 88
rect 258 87 260 96
rect 274 82 276 91
rect 284 82 286 91
rect 294 79 296 91
rect 301 79 303 91
rect 342 87 344 96
rect 358 82 360 91
rect 368 82 370 91
rect 378 79 380 91
rect 385 79 387 91
rect 412 85 414 91
rect 424 79 426 88
rect 431 79 433 88
rect 169 51 171 65
rect 180 45 182 65
rect 187 45 189 65
rect 207 45 209 59
rect 217 45 219 59
rect 227 52 229 62
rect 237 52 239 65
rect 273 51 275 57
rect 283 51 285 57
rect 293 51 295 57
<< ptransistor >>
rect 180 108 182 120
rect 190 108 192 118
rect 200 108 202 118
rect 266 109 268 136
rect 282 109 284 127
rect 292 109 294 127
rect 302 109 304 136
rect 350 109 352 136
rect 366 109 368 127
rect 376 109 378 127
rect 386 109 388 136
rect 412 108 414 120
rect 422 108 424 118
rect 432 108 434 118
rect 169 5 171 33
rect 179 5 181 33
rect 189 5 191 33
rect 207 8 209 33
rect 214 8 216 33
rect 224 17 226 30
rect 237 5 239 30
rect 273 6 275 24
rect 280 6 282 24
rect 293 15 295 27
<< polycontact >>
rect 191 124 195 128
rect 252 116 256 120
rect 181 100 185 104
rect 336 116 340 120
rect 289 101 293 105
rect 299 101 303 105
rect 423 124 427 128
rect 200 92 204 96
rect 268 95 272 99
rect 373 101 377 105
rect 383 101 387 105
rect 413 100 417 104
rect 352 95 356 99
rect 432 92 436 96
rect 168 37 172 41
rect 178 37 182 41
rect 188 37 192 41
rect 195 37 199 41
rect 214 37 218 41
rect 234 44 238 48
rect 228 34 232 38
rect 270 38 274 42
rect 282 38 286 42
rect 290 37 294 41
rect 280 30 284 34
<< ndcontact >>
rect 174 86 178 90
rect 252 91 256 95
rect 336 91 340 95
rect 203 83 207 87
rect 266 83 270 87
rect 278 86 282 90
rect 288 84 292 88
rect 185 74 189 78
rect 350 83 354 87
rect 362 86 366 90
rect 372 84 376 88
rect 306 74 310 78
rect 406 86 410 90
rect 435 83 439 87
rect 390 74 394 78
rect 417 74 421 78
rect 163 53 167 57
rect 174 60 178 64
rect 191 53 195 57
rect 201 53 205 57
rect 201 46 205 50
rect 211 46 215 50
rect 221 54 225 58
rect 231 57 235 61
rect 241 53 245 57
rect 267 52 271 56
rect 277 52 281 56
rect 287 52 291 56
rect 297 52 301 56
<< pdcontact >>
rect 174 109 178 113
rect 184 109 188 113
rect 194 109 198 113
rect 204 113 208 117
rect 260 110 264 114
rect 270 131 274 135
rect 270 124 274 128
rect 286 110 290 114
rect 296 117 300 121
rect 306 125 310 129
rect 344 110 348 114
rect 354 131 358 135
rect 354 124 358 128
rect 370 110 374 114
rect 380 117 384 121
rect 390 125 394 129
rect 406 109 410 113
rect 416 109 420 113
rect 426 109 430 113
rect 436 113 440 117
rect 163 28 167 32
rect 163 21 167 25
rect 173 13 177 17
rect 173 6 177 10
rect 183 21 187 25
rect 183 14 187 18
rect 195 13 199 17
rect 195 6 199 10
rect 218 25 222 29
rect 230 6 234 10
rect 241 25 245 29
rect 241 18 245 22
rect 267 14 271 18
rect 297 16 301 20
rect 285 7 289 11
<< m2contact >>
rect 197 124 201 128
rect 340 124 344 128
rect 173 96 177 100
rect 205 98 209 102
rect 242 98 246 102
rect 262 97 266 101
rect 309 97 313 101
rect 346 97 350 101
rect 429 124 433 128
rect 398 81 402 85
rect 437 99 441 103
rect 266 29 270 33
rect 257 21 261 25
<< psubstratepcontact >>
rect 175 74 179 78
rect 253 74 257 78
rect 337 74 341 78
rect 407 74 411 78
rect 268 64 272 68
rect 296 64 300 68
<< nsubstratencontact >>
rect 175 134 179 138
rect 189 134 193 138
rect 203 134 207 138
rect 286 134 290 138
rect 370 134 374 138
rect 407 134 411 138
rect 421 134 425 138
rect 435 134 439 138
rect 296 4 300 8
<< psubstratepdiff >>
rect 174 78 180 79
rect 174 74 175 78
rect 179 74 180 78
rect 174 73 180 74
rect 252 78 258 79
rect 252 74 253 78
rect 257 74 258 78
rect 252 73 258 74
rect 336 78 342 79
rect 336 74 337 78
rect 341 74 342 78
rect 336 73 342 74
rect 406 78 412 79
rect 406 74 407 78
rect 411 74 412 78
rect 406 73 412 74
rect 267 68 301 69
rect 267 64 268 68
rect 272 64 296 68
rect 300 64 301 68
rect 267 63 301 64
<< nsubstratendiff >>
rect 174 138 208 139
rect 174 134 175 138
rect 179 134 189 138
rect 193 134 203 138
rect 207 134 208 138
rect 285 138 291 139
rect 174 133 208 134
rect 285 134 286 138
rect 290 134 291 138
rect 369 138 375 139
rect 285 133 291 134
rect 369 134 370 138
rect 374 134 375 138
rect 406 138 440 139
rect 369 133 375 134
rect 406 134 407 138
rect 411 134 421 138
rect 425 134 435 138
rect 439 134 440 138
rect 406 133 440 134
rect 295 8 301 9
rect 295 4 296 8
rect 300 4 301 8
rect 295 3 301 4
<< pad >>
rect 175 53 179 57
<< labels >>
rlabel metal1 281 74 281 74 6 vss
rlabel metal1 281 138 281 138 6 vdd
rlabel metal1 365 74 365 74 6 vss
rlabel metal1 365 138 365 138 6 vdd
rlabel metal1 191 74 191 74 6 vss
rlabel metal1 191 138 191 138 6 vdd
rlabel metal1 423 138 423 138 6 vdd
rlabel metal1 423 74 423 74 6 vss
rlabel metal1 284 68 284 68 2 vss
rlabel metal1 284 4 284 4 2 vdd
rlabel metal1 196 106 196 106 1 co_n
rlabel metal1 183 86 183 86 1 co
rlabel metal1 407 102 407 102 1 c1
rlabel metal1 421 102 421 102 1 zc1_n
rlabel metal1 172 35 172 35 2 con
rlabel metal1 191 55 191 55 2 con
rlabel metal1 200 3 200 3 2 vdd
rlabel metal1 214 56 214 56 2 n2
rlabel metal1 203 52 203 52 2 n2
rlabel metal1 200 67 200 67 2 vss
rlabel metal1 230 30 230 30 2 con
rlabel metal1 220 29 220 29 2 son
rlabel polycontact 230 36 230 36 2 con
rlabel polycontact 269 98 269 98 1 a1
rlabel metal1 261 94 261 94 1 a1
rlabel metal1 253 122 253 122 1 b1
rlabel metal2 261 126 261 126 1 b1
rlabel metal1 254 100 254 100 1 b1n
rlabel ptransistor 293 111 293 111 1 a1n
rlabel metal1 309 106 309 106 1 x1
rlabel metal2 345 126 345 126 1 c0
rlabel metal1 393 106 393 106 1 s1
rlabel ntransistor 386 90 386 90 1 s1n
rlabel metal2 381 127 381 127 1 c0n
rlabel metal1 300 40 300 40 1 s2
rlabel metal1 292 36 292 36 1 s2n
rlabel polycontact 188 39 188 39 1 a0
rlabel metal2 188 31 188 31 1 b0
rlabel metal1 244 39 244 39 1 s0
<< end >>
